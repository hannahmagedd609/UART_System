module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX16M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX20M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX14M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX16M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX20M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY1X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1XLM (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MX2XLM (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFSRX2M (
	SN, 
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFSX1M (
	SN, 
	SI, 
	SE, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NAND3BXLM (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module INVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX2M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AO2B2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module BUFX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX4XLM (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSRX1M (
	SN, 
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND4XLM (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X1M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX12M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Fri Oct 25 20:28:13 2024
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_RST_N;
   wire FE_PHN6_RST_N;
   wire FE_PHN3_scan_rst;
   wire FE_PHN0_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC7_RST_N (
	.Y(FE_PHN7_RST_N),
	.A(FE_PHN6_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC6_RST_N (
	.Y(FE_PHN6_RST_N),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC3_scan_rst (
	.Y(FE_PHN3_scan_rst),
	.A(FE_PHN0_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_scan_rst (
	.Y(FE_PHN0_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN3_scan_rst),
	.A(FE_PHN7_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN5_scan_rst;
   wire FE_PHN2_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC5_scan_rst (
	.Y(FE_PHN5_scan_rst),
	.A(FE_PHN2_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_scan_rst (
	.Y(FE_PHN2_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN5_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN4_scan_rst;
   wire FE_PHN1_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC4_scan_rst (
	.Y(FE_PHN4_scan_rst),
	.A(FE_PHN1_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC1_scan_rst (
	.Y(FE_PHN1_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN4_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_1 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \RST_REG[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RST_REG_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\RST_REG[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RST_REG_reg[1]  (
	.SI(\RST_REG[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\RST_REG[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_0 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \RST_REG[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RST_REG_reg[1]  (
	.SI(\RST_REG[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\RST_REG[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RST_REG_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\RST_REG[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DATA_SYNC_BUS_WIDTH8_test_1 (
	unsync_bus, 
	bus_enable, 
	D_CLK, 
	RST, 
	sync_bus, 
	enable_pulse, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN3_O_RST2, 
	O_CLK1__L5_N7, 
	VDD, 
	VSS);
   input [7:0] unsync_bus;
   input bus_enable;
   input D_CLK;
   input RST;
   output [7:0] sync_bus;
   output enable_pulse;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN3_O_RST2;
   input O_CLK1__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n35;
   wire n18;
   wire n19;
   wire enable_flop;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n12;
   wire n17;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire [1:0] sync_flops;

   assign sync_bus[1] = n18 ;
   assign test_so = sync_flops[1] ;

   // Module instantiations
   INVXLM U3 (
	.Y(n10),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n35),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U5 (
	.Y(n12),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U6 (
	.Y(sync_bus[0]),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U7 (
	.Y(n17),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U11 (
	.Y(n1),
	.B(sync_flops[1]),
	.AN(enable_flop), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n6),
	.B1(n1),
	.B0(sync_bus[4]),
	.A1(n17),
	.A0(unsync_bus[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U13 (
	.Y(n2),
	.B1(n1),
	.B0(sync_bus[0]),
	.A1(n17),
	.A0(unsync_bus[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U14 (
	.Y(n3),
	.B1(n1),
	.B0(n35),
	.A1(n17),
	.A0(unsync_bus[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U15 (
	.Y(n4),
	.B1(n1),
	.B0(sync_bus[2]),
	.A1(n17),
	.A0(unsync_bus[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U16 (
	.Y(n7),
	.B1(n1),
	.B0(sync_bus[5]),
	.A1(n17),
	.A0(unsync_bus[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U17 (
	.Y(n5),
	.B1(n1),
	.B0(sync_bus[3]),
	.A1(n17),
	.A0(unsync_bus[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U18 (
	.Y(n8),
	.B1(n1),
	.B0(sync_bus[6]),
	.A1(n17),
	.A0(unsync_bus[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U19 (
	.Y(n9),
	.B1(n1),
	.B0(sync_bus[7]),
	.A1(n17),
	.A0(unsync_bus[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[7]  (
	.SI(sync_bus[6]),
	.SE(n25),
	.RN(RST),
	.Q(sync_bus[7]),
	.D(n9),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[6]  (
	.SI(sync_bus[5]),
	.SE(n24),
	.RN(RST),
	.Q(sync_bus[6]),
	.D(n8),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[5]  (
	.SI(sync_bus[4]),
	.SE(n30),
	.RN(RST),
	.Q(sync_bus[5]),
	.D(n7),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[3]  (
	.SI(sync_bus[2]),
	.SE(n30),
	.RN(FE_OFN3_O_RST2),
	.Q(sync_bus[3]),
	.D(n5),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_flops_reg[0]  (
	.SI(sync_bus[7]),
	.SE(n24),
	.RN(RST),
	.Q(sync_flops[0]),
	.D(bus_enable),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[2]  (
	.SI(n35),
	.SE(n29),
	.RN(FE_OFN3_O_RST2),
	.Q(sync_bus[2]),
	.D(n4),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_pulse_reg (
	.SI(enable_flop),
	.SE(n32),
	.RN(RST),
	.Q(enable_pulse),
	.D(n17),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_flops_reg[1]  (
	.SI(sync_flops[0]),
	.SE(n25),
	.RN(RST),
	.Q(sync_flops[1]),
	.D(sync_flops[0]),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_flop_reg (
	.SI(test_si),
	.SE(n31),
	.RN(RST),
	.Q(enable_flop),
	.D(sync_flops[1]),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[1]  (
	.SI(sync_bus[0]),
	.SE(n32),
	.RN(FE_OFN3_O_RST2),
	.Q(n18),
	.D(n3),
	.CK(D_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[0]  (
	.SI(enable_pulse),
	.SE(n31),
	.RN(RST),
	.Q(n19),
	.D(n2),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[4]  (
	.SI(sync_bus[3]),
	.SE(n29),
	.RN(FE_OFN3_O_RST2),
	.Q(sync_bus[4]),
	.D(n6),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U20 (
	.Y(n22),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U21 (
	.Y(n23),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U22 (
	.Y(n24),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U23 (
	.Y(n25),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U24 (
	.Y(n26),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U25 (
	.Y(n27),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U26 (
	.Y(n28),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U27 (
	.Y(n29),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U28 (
	.Y(n30),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U29 (
	.Y(n31),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U30 (
	.Y(n32),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ASYNC_FIFO_DATA_WIDTH8_ADD_WIDTH4_test_1 (
	W_CLK, 
	W_RST, 
	W_INC, 
	R_CLK, 
	R_RST, 
	R_INC, 
	WR_DATA, 
	FULL, 
	RD_DATA, 
	EMPTY, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN2_O_RST2, 
	FE_OFN3_O_RST2, 
	O_CLK3__L3_N3, 
	O_CLK1__L5_N5, 
	O_CLK1__L5_N6, 
	O_CLK1__L5_N7, 
	VDD, 
	VSS);
   input W_CLK;
   input W_RST;
   input W_INC;
   input R_CLK;
   input R_RST;
   input R_INC;
   input [7:0] WR_DATA;
   output FULL;
   output [7:0] RD_DATA;
   output EMPTY;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN2_O_RST2;
   input FE_OFN3_O_RST2;
   input O_CLK3__L3_N3;
   input O_CLK1__L5_N5;
   input O_CLK1__L5_N6;
   input O_CLK1__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n6;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire [2:0] waddr;
   wire [2:0] raddr;
   wire [3:0] wptr;
   wire [3:0] rq2_wptr;
   wire [3:0] rptr;
   wire [3:0] wq2_rptr;

   assign test_so2 = rptr[3] ;

   // Module instantiations
   DLY1X1M U9 (
	.Y(n10),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U10 (
	.Y(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U11 (
	.Y(n12),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U12 (
	.Y(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U13 (
	.Y(n14),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U14 (
	.Y(n15),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U15 (
	.Y(n16),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_MEM_CTRL_test_1 U0 (
	.w_data({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.W_CLK(W_CLK),
	.W_RST(W_RST),
	.w_addr({ waddr[2],
		waddr[1],
		waddr[0] }),
	.r_addr({ raddr[2],
		raddr[1],
		raddr[0] }),
	.winc(W_INC),
	.wfull(FULL),
	.r_data({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.test_si(test_si1),
	.test_so(n6),
	.test_se(n16),
	.FE_OFN2_O_RST2(FE_OFN2_O_RST2),
	.FE_OFN3_O_RST2(FE_OFN3_O_RST2),
	.O_CLK1__L5_N5(O_CLK1__L5_N5),
	.O_CLK1__L5_N6(O_CLK1__L5_N6),
	.O_CLK1__L5_N7(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_test_0 U1 (
	.in_ptr({ wptr[3],
		wptr[2],
		wptr[1],
		wptr[0] }),
	.CLK(R_CLK),
	.RST(R_RST),
	.out_ptr({ rq2_wptr[3],
		rq2_wptr[2],
		rq2_wptr[1],
		rq2_wptr[0] }),
	.test_si2(test_si2),
	.test_si1(n6),
	.test_so1(test_so1),
	.test_se(n13),
	.O_CLK3__L3_N3(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_test_1 U2 (
	.in_ptr({ rptr[3],
		rptr[2],
		rptr[1],
		rptr[0] }),
	.CLK(W_CLK),
	.RST(W_RST),
	.out_ptr({ wq2_rptr[3],
		wq2_rptr[2],
		wq2_rptr[1],
		wq2_rptr[0] }),
	.test_si(rq2_wptr[3]),
	.test_se(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_WR_test_1 U3 (
	.winc(W_INC),
	.wq2_rptr({ wq2_rptr[3],
		wq2_rptr[2],
		wq2_rptr[1],
		wq2_rptr[0] }),
	.W_CLK(W_CLK),
	.W_RST(W_RST),
	.wfull(FULL),
	.waddr({ waddr[2],
		waddr[1],
		waddr[0] }),
	.wptr({ wptr[3],
		wptr[2],
		wptr[1],
		wptr[0] }),
	.test_se(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_RD_test_1 U4 (
	.rinc(R_INC),
	.rq2_wptr({ rq2_wptr[3],
		rq2_wptr[2],
		rq2_wptr[1],
		rq2_wptr[0] }),
	.R_CLK(R_CLK),
	.R_RST(R_RST),
	.rempty(EMPTY),
	.raddr({ raddr[2],
		raddr[1],
		raddr[0] }),
	.rptr({ rptr[3],
		rptr[2],
		rptr[1],
		rptr[0] }),
	.test_si(wptr[3]),
	.test_se(n15),
	.O_CLK3__L3_N3(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_MEM_CTRL_test_1 (
	w_data, 
	W_CLK, 
	W_RST, 
	w_addr, 
	r_addr, 
	winc, 
	wfull, 
	r_data, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN2_O_RST2, 
	FE_OFN3_O_RST2, 
	O_CLK1__L5_N5, 
	O_CLK1__L5_N6, 
	O_CLK1__L5_N7, 
	VDD, 
	VSS);
   input [7:0] w_data;
   input W_CLK;
   input W_RST;
   input [2:0] w_addr;
   input [2:0] r_addr;
   input winc;
   input wfull;
   output [7:0] r_data;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN2_O_RST2;
   input FE_OFN3_O_RST2;
   input O_CLK1__L5_N5;
   input O_CLK1__L5_N6;
   input O_CLK1__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N10;
   wire N11;
   wire N12;
   wire \FIFO_Memory[0][7] ;
   wire \FIFO_Memory[0][6] ;
   wire \FIFO_Memory[0][5] ;
   wire \FIFO_Memory[0][4] ;
   wire \FIFO_Memory[0][3] ;
   wire \FIFO_Memory[0][2] ;
   wire \FIFO_Memory[0][1] ;
   wire \FIFO_Memory[0][0] ;
   wire \FIFO_Memory[1][7] ;
   wire \FIFO_Memory[1][6] ;
   wire \FIFO_Memory[1][5] ;
   wire \FIFO_Memory[1][4] ;
   wire \FIFO_Memory[1][3] ;
   wire \FIFO_Memory[1][2] ;
   wire \FIFO_Memory[1][1] ;
   wire \FIFO_Memory[1][0] ;
   wire \FIFO_Memory[2][7] ;
   wire \FIFO_Memory[2][6] ;
   wire \FIFO_Memory[2][5] ;
   wire \FIFO_Memory[2][4] ;
   wire \FIFO_Memory[2][3] ;
   wire \FIFO_Memory[2][2] ;
   wire \FIFO_Memory[2][1] ;
   wire \FIFO_Memory[2][0] ;
   wire \FIFO_Memory[3][7] ;
   wire \FIFO_Memory[3][6] ;
   wire \FIFO_Memory[3][5] ;
   wire \FIFO_Memory[3][4] ;
   wire \FIFO_Memory[3][3] ;
   wire \FIFO_Memory[3][2] ;
   wire \FIFO_Memory[3][1] ;
   wire \FIFO_Memory[3][0] ;
   wire \FIFO_Memory[4][7] ;
   wire \FIFO_Memory[4][6] ;
   wire \FIFO_Memory[4][5] ;
   wire \FIFO_Memory[4][4] ;
   wire \FIFO_Memory[4][3] ;
   wire \FIFO_Memory[4][2] ;
   wire \FIFO_Memory[4][1] ;
   wire \FIFO_Memory[4][0] ;
   wire \FIFO_Memory[5][7] ;
   wire \FIFO_Memory[5][6] ;
   wire \FIFO_Memory[5][5] ;
   wire \FIFO_Memory[5][4] ;
   wire \FIFO_Memory[5][3] ;
   wire \FIFO_Memory[5][2] ;
   wire \FIFO_Memory[5][1] ;
   wire \FIFO_Memory[5][0] ;
   wire \FIFO_Memory[6][7] ;
   wire \FIFO_Memory[6][6] ;
   wire \FIFO_Memory[6][5] ;
   wire \FIFO_Memory[6][4] ;
   wire \FIFO_Memory[6][3] ;
   wire \FIFO_Memory[6][2] ;
   wire \FIFO_Memory[6][1] ;
   wire \FIFO_Memory[6][0] ;
   wire \FIFO_Memory[7][7] ;
   wire \FIFO_Memory[7][6] ;
   wire \FIFO_Memory[7][5] ;
   wire \FIFO_Memory[7][4] ;
   wire \FIFO_Memory[7][3] ;
   wire \FIFO_Memory[7][2] ;
   wire \FIFO_Memory[7][1] ;
   wire \FIFO_Memory[7][0] ;
   wire n12;
   wire n16;
   wire n18;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n13;
   wire n14;
   wire n15;
   wire n17;
   wire n19;
   wire n20;
   wire n21;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n93;
   wire n94;
   wire n96;
   wire n97;
   wire n99;
   wire n101;
   wire n103;
   wire n105;
   wire n107;
   wire n109;
   wire n111;
   wire n113;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n177;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;

   assign N10 = r_addr[0] ;
   assign N11 = r_addr[1] ;
   assign N12 = r_addr[2] ;
   assign test_so = \FIFO_Memory[7][7]  ;

   // Module instantiations
   NOR2BX2M U2 (
	.Y(n18),
	.B(w_addr[2]),
	.AN(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n12),
	.B(n16),
	.A(w_addr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n131),
	.A(w_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n130),
	.A(w_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U13 (
	.Y(n99),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U15 (
	.Y(n107),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U18 (
	.Y(n16),
	.B(wfull),
	.AN(winc), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U19 (
	.Y(n105),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U21 (
	.Y(n103),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U23 (
	.Y(n101),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U25 (
	.Y(n1),
	.C(n18),
	.B(n131),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U26 (
	.Y(n2),
	.C(n12),
	.B(n131),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U27 (
	.Y(n109),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U29 (
	.Y(n111),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U31 (
	.Y(n113),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX4M U33 (
	.Y(n93),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U35 (
	.Y(n96),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U37 (
	.Y(n3),
	.C(n18),
	.B(n131),
	.A(w_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U38 (
	.Y(n54),
	.B1(n105),
	.B0(n129),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U39 (
	.Y(n55),
	.B1(n105),
	.B0(n122),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U40 (
	.Y(n56),
	.B1(n105),
	.B0(n123),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U41 (
	.Y(n57),
	.B1(n105),
	.B0(n124),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U42 (
	.Y(n58),
	.B1(n105),
	.B0(n125),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U43 (
	.Y(n59),
	.B1(n105),
	.B0(n126),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U44 (
	.Y(n60),
	.B1(n105),
	.B0(n127),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U45 (
	.Y(n61),
	.B1(n105),
	.B0(n128),
	.A1N(n105),
	.A0N(\FIFO_Memory[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U46 (
	.Y(n62),
	.B1(n103),
	.B0(n129),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U47 (
	.Y(n63),
	.B1(n103),
	.B0(n122),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U48 (
	.Y(n64),
	.B1(n103),
	.B0(n123),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U49 (
	.Y(n65),
	.B1(n103),
	.B0(n124),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U50 (
	.Y(n66),
	.B1(n103),
	.B0(n125),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U51 (
	.Y(n67),
	.B1(n103),
	.B0(n126),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U52 (
	.Y(n68),
	.B1(n103),
	.B0(n127),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U53 (
	.Y(n69),
	.B1(n103),
	.B0(n128),
	.A1N(n103),
	.A0N(\FIFO_Memory[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U54 (
	.Y(n70),
	.B1(n101),
	.B0(n129),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U55 (
	.Y(n71),
	.B1(n101),
	.B0(n122),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U56 (
	.Y(n72),
	.B1(n101),
	.B0(n123),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U57 (
	.Y(n73),
	.B1(n101),
	.B0(n124),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U58 (
	.Y(n74),
	.B1(n101),
	.B0(n125),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U59 (
	.Y(n75),
	.B1(n101),
	.B0(n126),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U60 (
	.Y(n76),
	.B1(n101),
	.B0(n127),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U61 (
	.Y(n77),
	.B1(n101),
	.B0(n128),
	.A1N(n101),
	.A0N(\FIFO_Memory[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U62 (
	.Y(n78),
	.B1(n99),
	.B0(n129),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U63 (
	.Y(n79),
	.B1(n99),
	.B0(n122),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U64 (
	.Y(n80),
	.B1(n99),
	.B0(n123),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U65 (
	.Y(n81),
	.B1(n99),
	.B0(n124),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U66 (
	.Y(n82),
	.B1(n99),
	.B0(n125),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U67 (
	.Y(n83),
	.B1(n99),
	.B0(n126),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U68 (
	.Y(n84),
	.B1(n99),
	.B0(n127),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U69 (
	.Y(n85),
	.B1(n99),
	.B0(n128),
	.A1N(n99),
	.A0N(\FIFO_Memory[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U70 (
	.Y(n4),
	.C(n18),
	.B(w_addr[0]),
	.A(w_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U71 (
	.Y(n5),
	.C(n18),
	.B(n130),
	.A(w_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U72 (
	.Y(n129),
	.A(w_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U73 (
	.Y(n122),
	.A(w_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U74 (
	.Y(n123),
	.A(w_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U75 (
	.Y(n124),
	.A(w_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U76 (
	.Y(n125),
	.A(w_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U77 (
	.Y(n126),
	.A(w_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U78 (
	.Y(n127),
	.A(w_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U79 (
	.Y(n128),
	.A(w_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U80 (
	.Y(n6),
	.C(w_addr[1]),
	.B(n12),
	.A(w_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U81 (
	.Y(n30),
	.B1(n111),
	.B0(n129),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U82 (
	.Y(n31),
	.B1(n111),
	.B0(n122),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U83 (
	.Y(n32),
	.B1(n111),
	.B0(n123),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n33),
	.B1(n111),
	.B0(n124),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n34),
	.B1(n111),
	.B0(n125),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n35),
	.B1(n111),
	.B0(n126),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n36),
	.B1(n111),
	.B0(n127),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n37),
	.B1(n111),
	.B0(n128),
	.A1N(n111),
	.A0N(\FIFO_Memory[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n38),
	.B1(n109),
	.B0(n129),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n39),
	.B1(n109),
	.B0(n122),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n40),
	.B1(n109),
	.B0(n123),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U92 (
	.Y(n41),
	.B1(n109),
	.B0(n124),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U93 (
	.Y(n42),
	.B1(n109),
	.B0(n125),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U94 (
	.Y(n43),
	.B1(n109),
	.B0(n126),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n44),
	.B1(n109),
	.B0(n127),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U96 (
	.Y(n45),
	.B1(n109),
	.B0(n128),
	.A1N(n109),
	.A0N(\FIFO_Memory[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U97 (
	.Y(n46),
	.B1(n107),
	.B0(n129),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U98 (
	.Y(n47),
	.B1(n107),
	.B0(n122),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U99 (
	.Y(n48),
	.B1(n107),
	.B0(n123),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n49),
	.B1(n107),
	.B0(n124),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n50),
	.B1(n107),
	.B0(n125),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n51),
	.B1(n107),
	.B0(n126),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n52),
	.B1(n107),
	.B0(n127),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n53),
	.B1(n107),
	.B0(n128),
	.A1N(n107),
	.A0N(\FIFO_Memory[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U105 (
	.Y(n22),
	.B1(n129),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U106 (
	.Y(n23),
	.B1(n122),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U107 (
	.Y(n24),
	.B1(n123),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U108 (
	.Y(n25),
	.B1(n124),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U109 (
	.Y(n26),
	.B1(n125),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U110 (
	.Y(n27),
	.B1(n126),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U111 (
	.Y(n28),
	.B1(n127),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U112 (
	.Y(n29),
	.B1(n128),
	.B0(n113),
	.A1N(n113),
	.A0N(\FIFO_Memory[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U113 (
	.Y(n7),
	.C(w_addr[0]),
	.B(n131),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U114 (
	.Y(n8),
	.C(w_addr[1]),
	.B(n130),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U115 (
	.Y(r_data[0]),
	.S0(n134),
	.B(n9),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U116 (
	.Y(n9),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][0] ),
	.C(\FIFO_Memory[6][0] ),
	.B(\FIFO_Memory[5][0] ),
	.A(\FIFO_Memory[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U117 (
	.Y(n10),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][0] ),
	.C(\FIFO_Memory[2][0] ),
	.B(\FIFO_Memory[1][0] ),
	.A(\FIFO_Memory[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U118 (
	.Y(r_data[1]),
	.S0(n177),
	.B(n11),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U119 (
	.Y(n11),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][1] ),
	.C(\FIFO_Memory[6][1] ),
	.B(\FIFO_Memory[5][1] ),
	.A(\FIFO_Memory[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U120 (
	.Y(n13),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][1] ),
	.C(\FIFO_Memory[2][1] ),
	.B(\FIFO_Memory[1][1] ),
	.A(\FIFO_Memory[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U121 (
	.Y(r_data[2]),
	.S0(n134),
	.B(n14),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U122 (
	.Y(n14),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][2] ),
	.C(\FIFO_Memory[6][2] ),
	.B(\FIFO_Memory[5][2] ),
	.A(\FIFO_Memory[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U123 (
	.Y(n15),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][2] ),
	.C(\FIFO_Memory[2][2] ),
	.B(\FIFO_Memory[1][2] ),
	.A(\FIFO_Memory[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U124 (
	.Y(r_data[3]),
	.S0(n134),
	.B(n17),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U125 (
	.Y(n17),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][3] ),
	.C(\FIFO_Memory[6][3] ),
	.B(\FIFO_Memory[5][3] ),
	.A(\FIFO_Memory[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U126 (
	.Y(n19),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][3] ),
	.C(\FIFO_Memory[2][3] ),
	.B(\FIFO_Memory[1][3] ),
	.A(\FIFO_Memory[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U127 (
	.Y(r_data[4]),
	.S0(n177),
	.B(n20),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U128 (
	.Y(n20),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][4] ),
	.C(\FIFO_Memory[6][4] ),
	.B(\FIFO_Memory[5][4] ),
	.A(\FIFO_Memory[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U129 (
	.Y(n21),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][4] ),
	.C(\FIFO_Memory[2][4] ),
	.B(\FIFO_Memory[1][4] ),
	.A(\FIFO_Memory[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U130 (
	.Y(r_data[5]),
	.S0(n134),
	.B(n86),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U131 (
	.Y(n86),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][5] ),
	.C(\FIFO_Memory[6][5] ),
	.B(\FIFO_Memory[5][5] ),
	.A(\FIFO_Memory[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U132 (
	.Y(n87),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][5] ),
	.C(\FIFO_Memory[2][5] ),
	.B(\FIFO_Memory[1][5] ),
	.A(\FIFO_Memory[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U133 (
	.Y(r_data[6]),
	.S0(n134),
	.B(n88),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U134 (
	.Y(n88),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][6] ),
	.C(\FIFO_Memory[6][6] ),
	.B(\FIFO_Memory[5][6] ),
	.A(\FIFO_Memory[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U135 (
	.Y(n89),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][6] ),
	.C(\FIFO_Memory[2][6] ),
	.B(\FIFO_Memory[1][6] ),
	.A(\FIFO_Memory[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U136 (
	.Y(r_data[7]),
	.S0(n177),
	.B(n90),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U137 (
	.Y(n90),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[7][7] ),
	.C(\FIFO_Memory[6][7] ),
	.B(\FIFO_Memory[5][7] ),
	.A(\FIFO_Memory[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U138 (
	.Y(n91),
	.S1(n96),
	.S0(n93),
	.D(\FIFO_Memory[3][7] ),
	.C(\FIFO_Memory[2][7] ),
	.B(\FIFO_Memory[1][7] ),
	.A(\FIFO_Memory[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U139 (
	.Y(n94),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U140 (
	.Y(n97),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][7]  (
	.SI(\FIFO_Memory[1][6] ),
	.SE(n184),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][7] ),
	.D(n77),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][6]  (
	.SI(\FIFO_Memory[1][5] ),
	.SE(n135),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][6] ),
	.D(n76),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][5]  (
	.SI(\FIFO_Memory[1][4] ),
	.SE(n183),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][5] ),
	.D(n75),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][4]  (
	.SI(\FIFO_Memory[1][3] ),
	.SE(n175),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][4] ),
	.D(n74),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][3]  (
	.SI(\FIFO_Memory[1][2] ),
	.SE(n160),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[1][3] ),
	.D(n73),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][2]  (
	.SI(\FIFO_Memory[1][1] ),
	.SE(n159),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][2] ),
	.D(n72),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][1]  (
	.SI(\FIFO_Memory[1][0] ),
	.SE(n172),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][1] ),
	.D(n71),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[1][0]  (
	.SI(\FIFO_Memory[0][7] ),
	.SE(n174),
	.RN(W_RST),
	.Q(\FIFO_Memory[1][0] ),
	.D(n70),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][1]  (
	.SI(\FIFO_Memory[2][0] ),
	.SE(n185),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][1] ),
	.D(n63),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][0]  (
	.SI(\FIFO_Memory[1][7] ),
	.SE(n136),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][0] ),
	.D(n62),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][7]  (
	.SI(\FIFO_Memory[0][6] ),
	.SE(n160),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][7] ),
	.D(n85),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][6]  (
	.SI(\FIFO_Memory[0][5] ),
	.SE(n159),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][6] ),
	.D(n84),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][5]  (
	.SI(\FIFO_Memory[0][4] ),
	.SE(n173),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][5] ),
	.D(n83),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][4]  (
	.SI(\FIFO_Memory[0][3] ),
	.SE(n175),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][4] ),
	.D(n82),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][3]  (
	.SI(\FIFO_Memory[0][2] ),
	.SE(n182),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][3] ),
	.D(n81),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][2]  (
	.SI(\FIFO_Memory[0][1] ),
	.SE(n181),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][2] ),
	.D(n80),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][1]  (
	.SI(\FIFO_Memory[0][0] ),
	.SE(n172),
	.RN(W_RST),
	.Q(\FIFO_Memory[0][1] ),
	.D(n79),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[0][0]  (
	.SI(test_si),
	.SE(n174),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[0][0] ),
	.D(n78),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][7]  (
	.SI(\FIFO_Memory[4][6] ),
	.SE(n196),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][7] ),
	.D(n53),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][6]  (
	.SI(\FIFO_Memory[4][5] ),
	.SE(n147),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][6] ),
	.D(n52),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][5]  (
	.SI(\FIFO_Memory[4][4] ),
	.SE(n195),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][5] ),
	.D(n51),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][4]  (
	.SI(\FIFO_Memory[4][3] ),
	.SE(n146),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][4] ),
	.D(n50),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][3]  (
	.SI(\FIFO_Memory[4][2] ),
	.SE(n194),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][3] ),
	.D(n49),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][2]  (
	.SI(\FIFO_Memory[4][1] ),
	.SE(n145),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][2] ),
	.D(n48),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][1]  (
	.SI(\FIFO_Memory[4][0] ),
	.SE(n193),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[4][1] ),
	.D(n47),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[4][0]  (
	.SI(\FIFO_Memory[3][7] ),
	.SE(n144),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[4][0] ),
	.D(n46),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][7]  (
	.SI(\FIFO_Memory[6][6] ),
	.SE(n204),
	.RN(W_RST),
	.Q(\FIFO_Memory[6][7] ),
	.D(n37),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][6]  (
	.SI(\FIFO_Memory[6][5] ),
	.SE(n155),
	.RN(W_RST),
	.Q(\FIFO_Memory[6][6] ),
	.D(n36),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][5]  (
	.SI(\FIFO_Memory[6][4] ),
	.SE(n203),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[6][5] ),
	.D(n35),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][4]  (
	.SI(\FIFO_Memory[6][3] ),
	.SE(n154),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[6][4] ),
	.D(n34),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][3]  (
	.SI(\FIFO_Memory[6][2] ),
	.SE(n202),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[6][3] ),
	.D(n33),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][2]  (
	.SI(\FIFO_Memory[6][1] ),
	.SE(n153),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[6][2] ),
	.D(n32),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][1]  (
	.SI(\FIFO_Memory[6][0] ),
	.SE(n201),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[6][1] ),
	.D(n31),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[6][0]  (
	.SI(\FIFO_Memory[5][7] ),
	.SE(n152),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[6][0] ),
	.D(n30),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][7]  (
	.SI(\FIFO_Memory[5][6] ),
	.SE(n200),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[5][7] ),
	.D(n45),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][6]  (
	.SI(\FIFO_Memory[5][5] ),
	.SE(n151),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[5][6] ),
	.D(n44),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][5]  (
	.SI(\FIFO_Memory[5][4] ),
	.SE(n199),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[5][5] ),
	.D(n43),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][4]  (
	.SI(\FIFO_Memory[5][3] ),
	.SE(n150),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[5][4] ),
	.D(n42),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][3]  (
	.SI(\FIFO_Memory[5][2] ),
	.SE(n198),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[5][3] ),
	.D(n41),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][2]  (
	.SI(\FIFO_Memory[5][1] ),
	.SE(n149),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[5][2] ),
	.D(n40),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][1]  (
	.SI(\FIFO_Memory[5][0] ),
	.SE(n197),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[5][1] ),
	.D(n39),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[5][0]  (
	.SI(\FIFO_Memory[4][7] ),
	.SE(n148),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[5][0] ),
	.D(n38),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][7]  (
	.SI(\FIFO_Memory[7][6] ),
	.SE(n161),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[7][7] ),
	.D(n29),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][6]  (
	.SI(\FIFO_Memory[7][5] ),
	.SE(n161),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[7][6] ),
	.D(n28),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][5]  (
	.SI(\FIFO_Memory[7][4] ),
	.SE(n207),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[7][5] ),
	.D(n27),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][4]  (
	.SI(\FIFO_Memory[7][3] ),
	.SE(n158),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[7][4] ),
	.D(n26),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][3]  (
	.SI(\FIFO_Memory[7][2] ),
	.SE(n206),
	.RN(FE_OFN3_O_RST2),
	.Q(\FIFO_Memory[7][3] ),
	.D(n25),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][2]  (
	.SI(\FIFO_Memory[7][1] ),
	.SE(n157),
	.RN(W_RST),
	.Q(\FIFO_Memory[7][2] ),
	.D(n24),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][1]  (
	.SI(\FIFO_Memory[7][0] ),
	.SE(n205),
	.RN(W_RST),
	.Q(\FIFO_Memory[7][1] ),
	.D(n23),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[7][0]  (
	.SI(\FIFO_Memory[6][7] ),
	.SE(n156),
	.RN(W_RST),
	.Q(\FIFO_Memory[7][0] ),
	.D(n22),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][7]  (
	.SI(\FIFO_Memory[3][6] ),
	.SE(n192),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][7] ),
	.D(n61),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][6]  (
	.SI(\FIFO_Memory[3][5] ),
	.SE(n143),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][6] ),
	.D(n60),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][5]  (
	.SI(\FIFO_Memory[3][4] ),
	.SE(n191),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][5] ),
	.D(n59),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][4]  (
	.SI(\FIFO_Memory[3][3] ),
	.SE(n142),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][4] ),
	.D(n58),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][3]  (
	.SI(\FIFO_Memory[3][2] ),
	.SE(n190),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][3] ),
	.D(n57),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][2]  (
	.SI(\FIFO_Memory[3][1] ),
	.SE(n141),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][2] ),
	.D(n56),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][1]  (
	.SI(\FIFO_Memory[3][0] ),
	.SE(n189),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][1] ),
	.D(n55),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[3][0]  (
	.SI(\FIFO_Memory[2][7] ),
	.SE(n140),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[3][0] ),
	.D(n54),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][7]  (
	.SI(\FIFO_Memory[2][6] ),
	.SE(n188),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][7] ),
	.D(n69),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][6]  (
	.SI(\FIFO_Memory[2][5] ),
	.SE(n139),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][6] ),
	.D(n68),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][5]  (
	.SI(\FIFO_Memory[2][4] ),
	.SE(n187),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][5] ),
	.D(n67),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][4]  (
	.SI(\FIFO_Memory[2][3] ),
	.SE(n138),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][4] ),
	.D(n66),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][3]  (
	.SI(\FIFO_Memory[2][2] ),
	.SE(n186),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][3] ),
	.D(n65),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FIFO_Memory_reg[2][2]  (
	.SI(\FIFO_Memory[2][1] ),
	.SE(n137),
	.RN(FE_OFN2_O_RST2),
	.Q(\FIFO_Memory[2][2] ),
	.D(n64),
	.CK(O_CLK1__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U141 (
	.Y(n134),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U142 (
	.Y(n135),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U143 (
	.Y(n136),
	.A(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U144 (
	.Y(n137),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U145 (
	.Y(n138),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U146 (
	.Y(n139),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U147 (
	.Y(n140),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U148 (
	.Y(n141),
	.A(n189), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U149 (
	.Y(n142),
	.A(n190), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U150 (
	.Y(n143),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U151 (
	.Y(n144),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U152 (
	.Y(n145),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U153 (
	.Y(n146),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U154 (
	.Y(n147),
	.A(n195), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U155 (
	.Y(n148),
	.A(n196), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U156 (
	.Y(n149),
	.A(n197), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U157 (
	.Y(n150),
	.A(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U158 (
	.Y(n151),
	.A(n199), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U159 (
	.Y(n152),
	.A(n200), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U160 (
	.Y(n153),
	.A(n201), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U161 (
	.Y(n154),
	.A(n202), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U162 (
	.Y(n155),
	.A(n203), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U163 (
	.Y(n156),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U164 (
	.Y(n157),
	.A(n205), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U165 (
	.Y(n158),
	.A(n206), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U166 (
	.Y(n159),
	.A(n181), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U167 (
	.Y(n160),
	.A(n182), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U168 (
	.Y(n161),
	.A(n207), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U177 (
	.Y(n170),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U178 (
	.Y(n171),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U179 (
	.Y(n172),
	.A(n180), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U180 (
	.Y(n173),
	.A(n180), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U181 (
	.Y(n174),
	.A(n179), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U182 (
	.Y(n175),
	.A(n179), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U184 (
	.Y(n177),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U186 (
	.Y(n179),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U187 (
	.Y(n180),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U188 (
	.Y(n181),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U189 (
	.Y(n182),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U190 (
	.Y(n183),
	.A(n173), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U191 (
	.Y(n184),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U192 (
	.Y(n185),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U193 (
	.Y(n186),
	.A(n137), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U194 (
	.Y(n187),
	.A(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U195 (
	.Y(n188),
	.A(n139), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U196 (
	.Y(n189),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U197 (
	.Y(n190),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U198 (
	.Y(n191),
	.A(n142), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U199 (
	.Y(n192),
	.A(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U200 (
	.Y(n193),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U201 (
	.Y(n194),
	.A(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U202 (
	.Y(n195),
	.A(n146), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U203 (
	.Y(n196),
	.A(n147), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U204 (
	.Y(n197),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U205 (
	.Y(n198),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U206 (
	.Y(n199),
	.A(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U207 (
	.Y(n200),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U208 (
	.Y(n201),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U209 (
	.Y(n202),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U210 (
	.Y(n203),
	.A(n154), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U211 (
	.Y(n204),
	.A(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U212 (
	.Y(n205),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U213 (
	.Y(n206),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U214 (
	.Y(n207),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_test_0 (
	in_ptr, 
	CLK, 
	RST, 
	out_ptr, 
	test_si2, 
	test_si1, 
	test_so1, 
	test_se, 
	O_CLK3__L3_N3, 
	VDD, 
	VSS);
   input [3:0] in_ptr;
   input CLK;
   input RST;
   output [3:0] out_ptr;
   input test_si2;
   input test_si1;
   output test_so1;
   input test_se;
   input O_CLK3__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \SYNC_reg[3][0] ;
   wire \SYNC_reg[2][0] ;
   wire \SYNC_reg[1][0] ;
   wire \SYNC_reg[0][0] ;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n3;

   // Module instantiations
   SDFFRQX2M \SYNC_reg_reg[3][1]  (
	.SI(test_si2),
	.SE(n10),
	.RN(RST),
	.Q(out_ptr[3]),
	.D(test_so1),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[2][1]  (
	.SI(\SYNC_reg[2][0] ),
	.SE(n7),
	.RN(RST),
	.Q(out_ptr[2]),
	.D(\SYNC_reg[2][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[1][1]  (
	.SI(\SYNC_reg[1][0] ),
	.SE(n8),
	.RN(RST),
	.Q(out_ptr[1]),
	.D(\SYNC_reg[1][0] ),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[0][1]  (
	.SI(\SYNC_reg[0][0] ),
	.SE(n12),
	.RN(RST),
	.Q(out_ptr[0]),
	.D(\SYNC_reg[0][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[3][0]  (
	.SI(out_ptr[2]),
	.SE(n8),
	.RN(RST),
	.Q(\SYNC_reg[3][0] ),
	.D(in_ptr[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[2][0]  (
	.SI(out_ptr[1]),
	.SE(n12),
	.RN(RST),
	.Q(\SYNC_reg[2][0] ),
	.D(in_ptr[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[1][0]  (
	.SI(out_ptr[0]),
	.SE(n7),
	.RN(RST),
	.Q(\SYNC_reg[1][0] ),
	.D(in_ptr[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[0][0]  (
	.SI(test_si1),
	.SE(n11),
	.RN(RST),
	.Q(\SYNC_reg[0][0] ),
	.D(in_ptr[0]),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U5 (
	.Y(n6),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U6 (
	.Y(n7),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U7 (
	.Y(n8),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U8 (
	.Y(n9),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U9 (
	.Y(n10),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U10 (
	.Y(n11),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U11 (
	.Y(n12),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U12 (
	.Y(n3),
	.A(\SYNC_reg[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M U13 (
	.Y(test_so1),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_test_1 (
	in_ptr, 
	CLK, 
	RST, 
	out_ptr, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [3:0] in_ptr;
   input CLK;
   input RST;
   output [3:0] out_ptr;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \SYNC_reg[3][0] ;
   wire \SYNC_reg[2][0] ;
   wire \SYNC_reg[1][0] ;
   wire \SYNC_reg[0][0] ;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;

   // Module instantiations
   SDFFRQX2M \SYNC_reg_reg[3][1]  (
	.SI(\SYNC_reg[3][0] ),
	.SE(n7),
	.RN(RST),
	.Q(out_ptr[3]),
	.D(\SYNC_reg[3][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[2][1]  (
	.SI(\SYNC_reg[2][0] ),
	.SE(n11),
	.RN(RST),
	.Q(out_ptr[2]),
	.D(\SYNC_reg[2][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[1][1]  (
	.SI(\SYNC_reg[1][0] ),
	.SE(n6),
	.RN(RST),
	.Q(out_ptr[1]),
	.D(\SYNC_reg[1][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[0][1]  (
	.SI(\SYNC_reg[0][0] ),
	.SE(n10),
	.RN(RST),
	.Q(out_ptr[0]),
	.D(\SYNC_reg[0][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[3][0]  (
	.SI(out_ptr[2]),
	.SE(n6),
	.RN(RST),
	.Q(\SYNC_reg[3][0] ),
	.D(in_ptr[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[2][0]  (
	.SI(out_ptr[1]),
	.SE(n7),
	.RN(RST),
	.Q(\SYNC_reg[2][0] ),
	.D(in_ptr[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[1][0]  (
	.SI(out_ptr[0]),
	.SE(n11),
	.RN(RST),
	.Q(\SYNC_reg[1][0] ),
	.D(in_ptr[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg_reg[0][0]  (
	.SI(test_si),
	.SE(n9),
	.RN(RST),
	.Q(\SYNC_reg[0][0] ),
	.D(in_ptr[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U5 (
	.Y(n5),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U6 (
	.Y(n6),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U7 (
	.Y(n7),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U8 (
	.Y(n8),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U9 (
	.Y(n9),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U10 (
	.Y(n10),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U11 (
	.Y(n11),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_WR_test_1 (
	winc, 
	wq2_rptr, 
	W_CLK, 
	W_RST, 
	wfull, 
	waddr, 
	wptr, 
	test_se, 
	VDD, 
	VSS);
   input winc;
   input [3:0] wq2_rptr;
   input W_CLK;
   input W_RST;
   output wfull;
   output [2:0] waddr;
   output [3:0] wptr;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n34;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n1;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n51;
   wire [2:0] wptr_reg;

   // Module instantiations
   CLKXOR2X2M U3 (
	.Y(wptr[0]),
	.B(wptr_reg[1]),
	.A(wptr_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U4 (
	.Y(wptr[1]),
	.B(wptr_reg[1]),
	.A(wptr_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U5 (
	.Y(n17),
	.D(wptr_reg[2]),
	.C(wptr[3]),
	.B(wptr_reg[1]),
	.A(wptr_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U6 (
	.Y(n1),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U7 (
	.Y(wptr[3]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U12 (
	.Y(wfull),
	.D(n21),
	.C(n20),
	.B(n19),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U13 (
	.Y(n15),
	.C(waddr[2]),
	.B(waddr[0]),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n31),
	.A(winc), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(n11),
	.B0(n17),
	.A1(n31),
	.A0(wfull), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U18 (
	.Y(n14),
	.B0(n15),
	.A1(n31),
	.A0(wfull), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U19 (
	.Y(n22),
	.B0(n9),
	.A2(n33),
	.A1(wptr_reg[2]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U20 (
	.Y(n9),
	.B0(wptr_reg[2]),
	.A1(n10),
	.A0(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n33),
	.A(wptr_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(wptr[2]),
	.B(wptr_reg[2]),
	.A(wptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n21),
	.B(wptr[3]),
	.A(wq2_rptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U24 (
	.Y(n18),
	.B(wq2_rptr[1]),
	.A(wptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U25 (
	.Y(n20),
	.B(wptr[2]),
	.A(wq2_rptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U26 (
	.Y(n8),
	.C(wptr_reg[0]),
	.B(n17),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U27 (
	.Y(n19),
	.B(wq2_rptr[0]),
	.A(wptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n29),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U29 (
	.Y(n16),
	.B1(wptr[3]),
	.B0(n17),
	.A2(wptr_reg[1]),
	.A1(wptr_reg[2]),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n30),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U31 (
	.Y(n25),
	.B(waddr[0]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(n27),
	.B(wptr_reg[0]),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U33 (
	.Y(n24),
	.B0(n13),
	.A1(n12),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U34 (
	.Y(n13),
	.B0(n32),
	.A1(waddr[0]),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U35 (
	.Y(n12),
	.C(waddr[0]),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U36 (
	.Y(n23),
	.B1(n8),
	.B0(wptr_reg[1]),
	.A1N(wptr_reg[1]),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U37 (
	.Y(n26),
	.B1(n12),
	.B0(n32),
	.A1N(waddr[2]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U38 (
	.Y(n10),
	.B(n11),
	.A(wptr_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n32),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \waddr_reg[2]  (
	.SI(n32),
	.SE(n40),
	.RN(W_RST),
	.Q(waddr[2]),
	.D(n26),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg_reg[0]  (
	.SI(waddr[2]),
	.SE(n37),
	.RN(W_RST),
	.Q(wptr_reg[0]),
	.D(n27),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg_reg[2]  (
	.SI(n33),
	.SE(n40),
	.RN(W_RST),
	.Q(wptr_reg[2]),
	.D(n22),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg_reg[3]  (
	.SI(wptr_reg[2]),
	.SE(n37),
	.RN(W_RST),
	.Q(n34),
	.D(n29),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg_reg[1]  (
	.SI(wptr_reg[0]),
	.SE(n39),
	.RN(W_RST),
	.Q(wptr_reg[1]),
	.D(n23),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \waddr_reg[0]  (
	.SI(wq2_rptr[3]),
	.SE(n38),
	.RN(W_RST),
	.Q(waddr[0]),
	.D(n25),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \waddr_reg[1]  (
	.SI(waddr[0]),
	.SE(n39),
	.RN(W_RST),
	.Q(waddr[1]),
	.D(n24),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U40 (
	.Y(n36),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U41 (
	.Y(n37),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U42 (
	.Y(n38),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U43 (
	.Y(n39),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U44 (
	.Y(n40),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U55 (
	.Y(n51),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_RD_test_1 (
	rinc, 
	rq2_wptr, 
	R_CLK, 
	R_RST, 
	rempty, 
	raddr, 
	rptr, 
	test_si, 
	test_se, 
	O_CLK3__L3_N3, 
	VDD, 
	VSS);
   input rinc;
   input [3:0] rq2_wptr;
   input R_CLK;
   input R_RST;
   output rempty;
   output [2:0] raddr;
   output [3:0] rptr;
   input test_si;
   input test_se;
   input O_CLK3__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n61;
   wire n62;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n30;
   wire n31;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n38;
   wire n40;
   wire n47;
   wire n58;
   wire [2:0] rptr_reg;

   // Module instantiations
   NAND3X2M U3 (
	.Y(n15),
	.C(n61),
	.B(raddr[0]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U6 (
	.Y(n11),
	.B0(n17),
	.A1(n7),
	.A0(rempty), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U7 (
	.Y(n14),
	.B0(n15),
	.A1(n7),
	.A0(rempty), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U8 (
	.Y(rptr[0]),
	.B(rptr_reg[1]),
	.A(rptr_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U9 (
	.Y(rptr[1]),
	.B(rptr_reg[1]),
	.A(rptr_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U10 (
	.Y(rptr[2]),
	.B(rptr_reg[2]),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U11 (
	.Y(rempty),
	.D(n21),
	.C(n20),
	.B(n19),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U12 (
	.Y(n20),
	.B(rq2_wptr[3]),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U13 (
	.Y(n19),
	.B(rq2_wptr[0]),
	.A(rptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U14 (
	.Y(n21),
	.B(rq2_wptr[2]),
	.A(rptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U15 (
	.Y(n18),
	.B(rq2_wptr[1]),
	.A(rptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U16 (
	.Y(n22),
	.B0(n9),
	.A2(n6),
	.A1(rptr_reg[2]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(n9),
	.B0(rptr_reg[2]),
	.A1(n10),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n6),
	.A(rptr_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n3),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U20 (
	.Y(n16),
	.B1(n62),
	.B0(n17),
	.A2(rptr_reg[1]),
	.A1(rptr_reg[2]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n4),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U22 (
	.Y(n17),
	.D(rptr_reg[2]),
	.C(n62),
	.B(rptr_reg[1]),
	.A(rptr_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U23 (
	.Y(n8),
	.C(rptr_reg[0]),
	.B(n17),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U24 (
	.Y(n25),
	.B(n40),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U25 (
	.Y(n27),
	.B(rptr_reg[0]),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U26 (
	.Y(n12),
	.C(n36),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U27 (
	.Y(n23),
	.B1(n8),
	.B0(rptr_reg[1]),
	.A1N(rptr_reg[1]),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U28 (
	.Y(n26),
	.B1(n5),
	.B0(n12),
	.A1N(n47),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U29 (
	.Y(n24),
	.B0(n13),
	.A1(n38),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U30 (
	.Y(n13),
	.B0(n5),
	.A1(n36),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U31 (
	.Y(n10),
	.B(n11),
	.A(rptr_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n7),
	.A(rinc), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \raddr_reg[0]  (
	.SI(test_si),
	.SE(n34),
	.RN(R_RST),
	.Q(raddr[0]),
	.D(n25),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rptr_reg_reg[3]  (
	.SI(rptr_reg[2]),
	.SE(n31),
	.RN(R_RST),
	.Q(n62),
	.D(n3),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rptr_reg_reg[0]  (
	.SI(n47),
	.SE(n35),
	.RN(R_RST),
	.Q(rptr_reg[0]),
	.D(n27),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rptr_reg_reg[2]  (
	.SI(n6),
	.SE(n35),
	.RN(R_RST),
	.Q(rptr_reg[2]),
	.D(n22),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rptr_reg_reg[1]  (
	.SI(rptr_reg[0]),
	.SE(n31),
	.RN(R_RST),
	.Q(rptr_reg[1]),
	.D(n23),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \raddr_reg[1]  (
	.SI(n40),
	.SE(n33),
	.RN(R_RST),
	.QN(n5),
	.Q(raddr[1]),
	.D(n24),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U33 (
	.Y(n30),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U34 (
	.Y(n31),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U36 (
	.Y(n33),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U37 (
	.Y(n34),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U38 (
	.Y(n35),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U39 (
	.Y(n36),
	.A(raddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U41 (
	.Y(n38),
	.A(raddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U43 (
	.Y(n40),
	.A(raddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U45 (
	.Y(rptr[3]),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U50 (
	.Y(n47),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U60 (
	.Y(raddr[2]),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \raddr_reg[2]  (
	.SI(n5),
	.SE(n33),
	.RN(R_RST),
	.QN(n58),
	.Q(n61),
	.D(n26),
	.CK(O_CLK3__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GEN_test_1 (
	CLK, 
	RST, 
	LVL_SIG, 
	PULSE_SIG, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input LVL_SIG;
   output PULSE_SIG;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire pulse_flop;
   wire prev_flop;

   assign test_so = pulse_flop ;

   // Module instantiations
   NOR2BX2M U3 (
	.Y(PULSE_SIG),
	.B(pulse_flop),
	.AN(prev_flop), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M pulse_flop_reg (
	.SI(prev_flop),
	.SE(test_se),
	.RN(RST),
	.Q(pulse_flop),
	.D(prev_flop),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M prev_flop_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(prev_flop),
	.D(LVL_SIG),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_width8_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	O_CLK2__L13_N0, 
	O_CLK2__L7_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input O_CLK2__L13_N0;
   input O_CLK2__L7_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN11_n44;
   wire FE_PHN10_n44;
   wire output_clk__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire N0;
   wire output_clk;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire n16;
   wire n17;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n73;
   wire [7:0] cyc_counter;

   assign N22 = i_div_ratio[1] ;
   assign N23 = i_div_ratio[2] ;
   assign N24 = i_div_ratio[3] ;
   assign N25 = i_div_ratio[4] ;
   assign N26 = i_div_ratio[5] ;
   assign N27 = i_div_ratio[6] ;
   assign N28 = i_div_ratio[7] ;

   // Module instantiations
   DLY4X1M FE_PHC11_n44 (
	.Y(FE_PHN10_n44),
	.A(FE_PHN11_n44), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC10_n44 (
	.Y(n44),
	.A(FE_PHN10_n44), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M output_clk__Exclude_0 (
	.Y(output_clk__Exclude_0_NET),
	.A(output_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U3 (
	.Y(n31),
	.D(n35),
	.C(n34),
	.B(n33),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U4 (
	.Y(n21),
	.D(n24),
	.C(n15),
	.B(n23),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U5 (
	.Y(n22),
	.C(N0),
	.B(n73),
	.AN(cyc_counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U6 (
	.Y(N17),
	.C(n7),
	.B(n56),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U7 (
	.Y(n9),
	.C(n15),
	.B(n13),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U8 (
	.Y(n13),
	.D(n31),
	.C(n30),
	.B(n29),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U9 (
	.Y(n30),
	.C(n38),
	.B(n37),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U10 (
	.Y(n11),
	.D(n21),
	.C(n20),
	.B(n19),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U11 (
	.Y(n20),
	.C(n27),
	.B(n26),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U12 (
	.Y(n37),
	.B0(HTIE_LTIEHI_NET),
	.A1(n40),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U13 (
	.Y(n7),
	.B(n53),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U14 (
	.Y(n6),
	.B(n55),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U15 (
	.Y(n5),
	.B(n51),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1XLM U16 (
	.Y(N12),
	.B0(n5),
	.A1N(n51),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U20 (
	.Y(n12),
	.C0(n14),
	.B0(n11),
	.A1(n13),
	.A0(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U21 (
	.Y(n4),
	.B(n58),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U22 (
	.Y(o_div_clk),
	.S0(N0),
	.B(output_clk),
	.A(O_CLK2__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U23 (
	.Y(N10),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U24 (
	.Y(N11),
	.B0(n4),
	.A1N(n49),
	.A0N(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U25 (
	.Y(N13),
	.B0(n6),
	.A1N(n55),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U26 (
	.Y(N14),
	.B0(n7),
	.A1N(n53),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U27 (
	.Y(N15),
	.B(n7),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U28 (
	.Y(n8),
	.B0(n57),
	.A1(n7),
	.A0(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U29 (
	.Y(N16),
	.B(n8),
	.AN(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U30 (
	.Y(n17),
	.B0(n11),
	.A1(n73),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U31 (
	.Y(n16),
	.B(output_clk__Exclude_0_NET),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U32 (
	.Y(N50),
	.B(n12),
	.AN(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U33 (
	.Y(N49),
	.B(n12),
	.AN(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U34 (
	.Y(N48),
	.B(n12),
	.AN(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U35 (
	.Y(N47),
	.B(n12),
	.AN(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U36 (
	.Y(N46),
	.B(n12),
	.AN(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U37 (
	.Y(N45),
	.B(n12),
	.AN(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U38 (
	.Y(N44),
	.B(n12),
	.AN(N35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U39 (
	.Y(N43),
	.B(n12),
	.AN(N34), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U40 (
	.Y(n14),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(n24),
	.B(n48),
	.A(cyc_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U42 (
	.Y(n15),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n23),
	.B(n58),
	.A(cyc_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U44 (
	.Y(n27),
	.B(n50),
	.A(cyc_counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U45 (
	.Y(n26),
	.B(n52),
	.A(cyc_counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n25),
	.B(n54),
	.A(cyc_counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U47 (
	.Y(n19),
	.B(cyc_counter[5]),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U48 (
	.Y(n18),
	.B(cyc_counter[6]),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n35),
	.B(N16),
	.A(cyc_counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n34),
	.B(N15),
	.A(cyc_counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n33),
	.B(N14),
	.A(cyc_counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n32),
	.B(N13),
	.A(cyc_counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n38),
	.B(N11),
	.A(cyc_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n36),
	.B(cyc_counter[0]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n29),
	.B(N12),
	.A(cyc_counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U56 (
	.Y(n28),
	.B(N17),
	.A(cyc_counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U57 (
	.Y(N0),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X1M U58 (
	.Y(n40),
	.C(n45),
	.B(n50),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U59 (
	.Y(n39),
	.D(n57),
	.C(n61),
	.B(n52),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[7]  (
	.SI(cyc_counter[6]),
	.SE(n46),
	.RN(i_rst_n),
	.Q(cyc_counter[7]),
	.D(N50),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[2]  (
	.SI(cyc_counter[1]),
	.SE(n69),
	.RN(i_rst_n),
	.Q(cyc_counter[2]),
	.D(N45),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[6]  (
	.SI(cyc_counter[5]),
	.SE(n47),
	.RN(i_rst_n),
	.Q(cyc_counter[6]),
	.D(N49),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[5]  (
	.SI(cyc_counter[4]),
	.SE(n69),
	.RN(i_rst_n),
	.Q(cyc_counter[5]),
	.D(N48),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[4]  (
	.SI(cyc_counter[3]),
	.SE(n46),
	.RN(i_rst_n),
	.Q(cyc_counter[4]),
	.D(N47),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[3]  (
	.SI(cyc_counter[2]),
	.SE(n47),
	.RN(i_rst_n),
	.Q(cyc_counter[3]),
	.D(N46),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[1]  (
	.SI(cyc_counter[0]),
	.SE(n67),
	.RN(i_rst_n),
	.Q(cyc_counter[1]),
	.D(N44),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cyc_counter_reg[0]  (
	.SI(test_si),
	.SE(n68),
	.RN(i_rst_n),
	.Q(cyc_counter[0]),
	.D(N43),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U60 (
	.Y(n45),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U61 (
	.Y(n46),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U62 (
	.Y(n47),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U63 (
	.Y(n48),
	.A(N23), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U64 (
	.Y(n49),
	.A(N23), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U65 (
	.Y(n50),
	.A(N24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U66 (
	.Y(n51),
	.A(N24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U67 (
	.Y(n52),
	.A(N26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U68 (
	.Y(n53),
	.A(N26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U69 (
	.Y(n54),
	.A(N25), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U70 (
	.Y(n55),
	.A(N25), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U71 (
	.Y(n56),
	.A(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U72 (
	.Y(n57),
	.A(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U73 (
	.Y(n58),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U74 (
	.Y(n59),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U76 (
	.Y(n61),
	.A(N27), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U77 (
	.Y(n62),
	.A(N27), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U78 (
	.Y(n63),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U79 (
	.Y(n64),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U80 (
	.Y(n65),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U81 (
	.Y(n66),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U82 (
	.Y(n67),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U83 (
	.Y(n68),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U84 (
	.Y(n69),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_width8_DW01_inc_0 add_57 (
	.A({ cyc_counter[7],
		cyc_counter[6],
		cyc_counter[5],
		cyc_counter[4],
		cyc_counter[3],
		cyc_counter[2],
		cyc_counter[1],
		cyc_counter[0] }),
	.SUM({ N41,
		N40,
		N39,
		N38,
		N37,
		N36,
		N35,
		N34 }), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M x_flag_reg (
	.SN(HTIE_LTIEHI_NET),
	.SI(n44),
	.SE(n66),
	.RN(i_rst_n),
	.QN(n73),
	.Q(test_so),
	.D(n17),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M output_clk_reg (
	.SN(HTIE_LTIEHI_NET),
	.SI(cyc_counter[7]),
	.SE(n66),
	.RN(i_rst_n),
	.QN(FE_PHN11_n44),
	.Q(output_clk),
	.D(n16),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_width8_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Pres_MUX_WIDTH4_PRE_WD6 (
	Prescale, 
	div_ratio, 
	VDD, 
	VSS);
   input [5:0] Prescale;
   output [3:0] div_ratio;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n29;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n1;
   wire n2;
   wire n3;
   wire n21;
   wire n26;

   // Module instantiations
   NOR3X2M U6 (
	.Y(div_ratio[1]),
	.C(Prescale[0]),
	.B(Prescale[1]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U3 (
	.Y(n8),
	.D(n2),
	.C(Prescale[3]),
	.B(Prescale[4]),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U4 (
	.Y(n3),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U5 (
	.Y(div_ratio[2]),
	.C(Prescale[0]),
	.B(Prescale[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U7 (
	.Y(n7),
	.D(n1),
	.C(n2),
	.B(Prescale[4]),
	.AN(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U8 (
	.Y(n6),
	.D(n1),
	.C(n2),
	.B(Prescale[3]),
	.AN(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U10 (
	.Y(n5),
	.C(Prescale[2]),
	.B(n3),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U11 (
	.Y(div_ratio[0]),
	.C0(n3),
	.B0(n21),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U12 (
	.Y(n9),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n2),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n1),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U25 (
	.Y(n21),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U28 (
	.Y(div_ratio[3]),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U31 (
	.Y(n29),
	.D(Prescale[4]),
	.C(Prescale[5]),
	.B(Prescale[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U32 (
	.Y(n26),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_width4_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	O_CLK2__L13_N0, 
	O_CLK2__L7_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [3:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input O_CLK2__L13_N0;
   input O_CLK2__L7_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN9_n35;
   wire FE_PHN8_n35;
   wire output_clk__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire output_clk;
   wire x_flag;
   wire N18;
   wire N19;
   wire N20;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n1;
   wire n2;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n10;
   wire n13;
   wire n14;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n76;
   wire [3:0] cyc_counter;

   assign N18 = i_div_ratio[1] ;
   assign N19 = i_div_ratio[2] ;
   assign N20 = i_div_ratio[3] ;
   assign test_so = n41 ;

   // Module instantiations
   DLY4X1M FE_PHC9_n35 (
	.Y(FE_PHN8_n35),
	.A(FE_PHN9_n35), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC8_n35 (
	.Y(n35),
	.A(FE_PHN8_n35), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M output_clk__Exclude_0 (
	.Y(output_clk__Exclude_0_NET),
	.A(output_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U14 (
	.Y(n15),
	.C0(n17),
	.B0(n6),
	.A1(n22),
	.A0(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U3 (
	.Y(n27),
	.B0(HTIE_LTIEHI_NET),
	.A2(N19),
	.A1(n37),
	.A0(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U4 (
	.Y(n26),
	.D(n7),
	.C(n2),
	.B(cyc_counter[3]),
	.A(x_flag), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n1),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U6 (
	.Y(n2),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U7 (
	.Y(N34),
	.B1(n10),
	.B0(n19),
	.A2(n76),
	.A1(cyc_counter[3]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U8 (
	.Y(n21),
	.B(cyc_counter[1]),
	.A(cyc_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U9 (
	.Y(n23),
	.B(cyc_counter[1]),
	.A(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U10 (
	.Y(n18),
	.C(n5),
	.B(cyc_counter[0]),
	.A(cyc_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U11 (
	.Y(N31),
	.B(cyc_counter[0]),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U12 (
	.Y(n28),
	.C(N18),
	.B(N19),
	.A(cyc_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n6),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(n16),
	.C(n7),
	.B(n22),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(n31),
	.B(n32),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(n32),
	.B0(n37),
	.A1(N19),
	.A0(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(n24),
	.B(n76),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U19 (
	.Y(n34),
	.B0(n17),
	.A1(n41),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n7),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U23 (
	.Y(n19),
	.B(n76),
	.AN(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U24 (
	.Y(n20),
	.B0(N31),
	.A1N(n15),
	.A0N(cyc_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U25 (
	.Y(N33),
	.B1(n18),
	.B0(cyc_counter[2]),
	.A1(n76),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U26 (
	.Y(n33),
	.B(output_clk__Exclude_0_NET),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U27 (
	.Y(n22),
	.D(n30),
	.C(n29),
	.B(n28),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U28 (
	.Y(n30),
	.B(N18),
	.A(cyc_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(n29),
	.B(cyc_counter[3]),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n5),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U31 (
	.Y(n17),
	.D(n26),
	.C(n25),
	.B(n24),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(n25),
	.B(cyc_counter[0]),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(N32),
	.B(n15),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U34 (
	.Y(o_div_clk),
	.S0(n1),
	.B(output_clk),
	.A(O_CLK2__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U35 (
	.Y(n36),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U36 (
	.Y(n37),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U37 (
	.Y(n38),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U38 (
	.Y(n39),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U39 (
	.Y(n40),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U75 (
	.Y(n76),
	.A(cyc_counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M x_flag_reg (
	.SN(HTIE_LTIEHI_NET),
	.SI(n35),
	.SE(n40),
	.RN(i_rst_n),
	.QN(n41),
	.Q(x_flag),
	.D(n34),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M output_clk_reg (
	.SN(HTIE_LTIEHI_NET),
	.SI(n10),
	.SE(n39),
	.RN(i_rst_n),
	.QN(FE_PHN9_n35),
	.Q(output_clk),
	.D(n33),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M \cyc_counter_reg[0]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(test_si),
	.SE(n38),
	.RN(i_rst_n),
	.QN(n14),
	.Q(cyc_counter[0]),
	.D(N31),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M \cyc_counter_reg[1]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(n14),
	.SE(n39),
	.RN(i_rst_n),
	.QN(n13),
	.Q(cyc_counter[1]),
	.D(N32),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M \cyc_counter_reg[2]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(n13),
	.SE(n40),
	.RN(i_rst_n),
	.QN(n9),
	.Q(cyc_counter[2]),
	.D(N33),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M \cyc_counter_reg[3]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(cyc_counter[2]),
	.SE(n38),
	.RN(i_rst_n),
	.QN(n10),
	.Q(cyc_counter[3]),
	.D(N34),
	.CK(O_CLK2__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_DATA_WIDTH8_test_1 (
	RST, 
	TX_CLK, 
	RX_CLK, 
	RX_IN_S, 
	RX_OUT_P, 
	RX_OUT_V, 
	TX_IN_P, 
	TX_IN_V, 
	TX_OUT_S, 
	TX_OUT_V, 
	Prescale, 
	parity_enable, 
	parity_type, 
	parity_error, 
	framing_error, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	O_CLK4__L3_N1, 
	O_CLK3__L3_N2, 
	VDD, 
	VSS);
   input RST;
   input TX_CLK;
   input RX_CLK;
   input RX_IN_S;
   output [7:0] RX_OUT_P;
   output RX_OUT_V;
   input [7:0] TX_IN_P;
   input TX_IN_V;
   output TX_OUT_S;
   output TX_OUT_V;
   input [5:0] Prescale;
   input parity_enable;
   input parity_type;
   output parity_error;
   output framing_error;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input O_CLK4__L3_N1;
   input O_CLK3__L3_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN4_O_RST3;
   wire n5;
   wire n9;

   // Module instantiations
   BUFX4M FE_OFC4_O_RST3 (
	.Y(FE_OFN4_O_RST3),
	.A(RST), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U3 (
	.Y(n9),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_TOP_test_1 U0_UART_TX (
	.P_DATA_M({ TX_IN_P[7],
		TX_IN_P[6],
		TX_IN_P[5],
		TX_IN_P[4],
		TX_IN_P[3],
		TX_IN_P[2],
		TX_IN_P[1],
		TX_IN_P[0] }),
	.Data_Valid_M(TX_IN_V),
	.PAR_EN_M(parity_enable),
	.PAR_TYPE_M(parity_type),
	.CLK_M(TX_CLK),
	.RST_M(RST),
	.TX_OUT_M(TX_OUT_S),
	.Busy_M(TX_OUT_V),
	.test_si(test_si1),
	.test_so(n5),
	.test_se(n9),
	.FE_OFN4_O_RST3(FE_OFN4_O_RST3),
	.O_CLK3__L3_N2(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_RX_test_1 U1_UART_RX (
	.CLK(RX_CLK),
	.RST(RST),
	.RX_IN(RX_IN_S),
	.parity_enable(parity_enable),
	.parity_type(parity_type),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.P_DATA({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.data_valid(RX_OUT_V),
	.parity_error(parity_error),
	.framing_error(framing_error),
	.test_si2(test_si2),
	.test_si1(n5),
	.test_so2(test_so2),
	.test_so1(test_so1),
	.test_se(n9),
	.FE_OFN4_O_RST3(FE_OFN4_O_RST3),
	.O_CLK4__L3_N1(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_TOP_test_1 (
	P_DATA_M, 
	Data_Valid_M, 
	PAR_EN_M, 
	PAR_TYPE_M, 
	CLK_M, 
	RST_M, 
	TX_OUT_M, 
	Busy_M, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_O_RST3, 
	O_CLK3__L3_N2, 
	VDD, 
	VSS);
   input [7:0] P_DATA_M;
   input Data_Valid_M;
   input PAR_EN_M;
   input PAR_TYPE_M;
   input CLK_M;
   input RST_M;
   output TX_OUT_M;
   output Busy_M;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_O_RST3;
   input O_CLK3__L3_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire ser_en_M;
   wire ser_data_M;
   wire ser_done_M;
   wire par_bit_M;
   wire n5;
   wire n8;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire [1:0] mux_sel_M;

   // Module instantiations
   DLY1X1M U4 (
	.Y(n8),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U8 (
	.Y(n12),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U9 (
	.Y(n13),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U10 (
	.Y(n14),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U11 (
	.Y(n15),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_Serial_test_1 Serial_DUT (
	.P_DATA({ P_DATA_M[7],
		P_DATA_M[6],
		P_DATA_M[5],
		P_DATA_M[4],
		P_DATA_M[3],
		P_DATA_M[2],
		P_DATA_M[1],
		P_DATA_M[0] }),
	.Data_Valid(Data_Valid_M),
	.ser_en(ser_en_M),
	.CLK(CLK_M),
	.RST(FE_OFN4_O_RST3),
	.Busy(Busy_M),
	.ser_done(ser_done_M),
	.ser_data(ser_data_M),
	.test_si(par_bit_M),
	.test_so(test_so),
	.test_se(n15),
	.O_CLK3__L3_N2(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_T_FSM_test_1 FSM_DUT (
	.Data_Valid(Data_Valid_M),
	.PAR_EN(PAR_EN_M),
	.ser_done(ser_done_M),
	.CLK(CLK_M),
	.RST(RST_M),
	.mux_sel({ mux_sel_M[1],
		mux_sel_M[0] }),
	.Busy(Busy_M),
	.ser_en(ser_en_M),
	.test_si(test_si),
	.test_so(n5),
	.test_se(n14),
	.FE_OFN4_O_RST3(FE_OFN4_O_RST3),
	.O_CLK3__L3_N2(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_Parity_calc_test_1 Parity_calc_DUT (
	.P_DATA({ P_DATA_M[7],
		P_DATA_M[6],
		P_DATA_M[5],
		P_DATA_M[4],
		P_DATA_M[3],
		P_DATA_M[2],
		P_DATA_M[1],
		P_DATA_M[0] }),
	.Data_Valid(Data_Valid_M),
	.PAR_TYPE(PAR_TYPE_M),
	.PAR_EN(PAR_EN_M),
	.CLK(CLK_M),
	.RST(RST_M),
	.Busy(Busy_M),
	.par_bit(par_bit_M),
	.test_si(TX_OUT_M),
	.test_se(n13),
	.FE_OFN4_O_RST3(FE_OFN4_O_RST3), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_MUX_test_1 MUX_DUT (
	.mux_sel({ mux_sel_M[1],
		mux_sel_M[0] }),
	.start_bit(1'b0),
	.stop_bit(1'b0),
	.ser_data(ser_data_M),
	.par_bit(par_bit_M),
	.CLK(CLK_M),
	.RST(RST_M),
	.TX_OUT(TX_OUT_M),
	.test_si(n5),
	.test_se(n14), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_Serial_test_1 (
	P_DATA, 
	Data_Valid, 
	ser_en, 
	CLK, 
	RST, 
	Busy, 
	ser_done, 
	ser_data, 
	test_si, 
	test_so, 
	test_se, 
	O_CLK3__L3_N2, 
	VDD, 
	VSS);
   input [7:0] P_DATA;
   input Data_Valid;
   input ser_en;
   input CLK;
   input RST;
   input Busy;
   output ser_done;
   output ser_data;
   input test_si;
   output test_so;
   input test_se;
   input O_CLK3__L3_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n6;
   wire n7;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n1;
   wire n2;
   wire n8;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire [2:0] P_Counter;
   wire [7:1] Temp_Reg;

   // Module instantiations
   NAND2X2M U3 (
	.Y(n1),
	.B(n11),
	.A(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n8),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U8 (
	.Y(n6),
	.B(n2),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U9 (
	.Y(n2),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U10 (
	.Y(n12),
	.B0(n6),
	.A1(n33),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U11 (
	.Y(n32),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U12 (
	.Y(n21),
	.B1(n35),
	.B0(n10),
	.A2(n34),
	.A1(P_Counter[2]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U13 (
	.Y(n10),
	.B0N(n12),
	.A1(n11),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U14 (
	.Y(n23),
	.B1(n8),
	.B0(n33),
	.A2(n32),
	.A1(P_Counter[0]),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U15 (
	.Y(n11),
	.B(Data_Valid),
	.AN(Busy), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U16 (
	.Y(n22),
	.B1(P_Counter[1]),
	.B0(n9),
	.A1(n34),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U17 (
	.Y(n9),
	.C(P_Counter[0]),
	.B(n11),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U18 (
	.Y(n24),
	.B0(n13),
	.A1N(n6),
	.A0N(ser_data), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U19 (
	.Y(n13),
	.B1(n32),
	.B0(P_DATA[0]),
	.A1(n2),
	.A0(Temp_Reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U20 (
	.Y(n31),
	.B0(n19),
	.A1N(Temp_Reg[1]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U21 (
	.Y(n19),
	.B1(n32),
	.B0(P_DATA[1]),
	.A1(n2),
	.A0(Temp_Reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U22 (
	.Y(n30),
	.B0(n18),
	.A1N(Temp_Reg[2]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U23 (
	.Y(n18),
	.B1(n32),
	.B0(P_DATA[2]),
	.A1(n2),
	.A0(Temp_Reg[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U24 (
	.Y(n29),
	.B0(n17),
	.A1N(Temp_Reg[3]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U25 (
	.Y(n17),
	.B1(n32),
	.B0(P_DATA[3]),
	.A1(n2),
	.A0(Temp_Reg[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U26 (
	.Y(n28),
	.B0(n16),
	.A1N(Temp_Reg[4]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U27 (
	.Y(n16),
	.B1(n32),
	.B0(P_DATA[4]),
	.A1(n2),
	.A0(Temp_Reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U28 (
	.Y(n27),
	.B0(n15),
	.A1N(Temp_Reg[5]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U29 (
	.Y(n15),
	.B1(n32),
	.B0(P_DATA[5]),
	.A1(n2),
	.A0(Temp_Reg[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U30 (
	.Y(n26),
	.B0(n14),
	.A1N(Temp_Reg[6]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U31 (
	.Y(n14),
	.B1(n32),
	.B0(P_DATA[6]),
	.A1(n2),
	.A0(Temp_Reg[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U32 (
	.Y(n20),
	.B0(n7),
	.A1N(n49),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U33 (
	.Y(n7),
	.D(P_Counter[0]),
	.C(n2),
	.B(P_Counter[1]),
	.A(P_Counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U34 (
	.Y(n25),
	.B1(n32),
	.B0(P_DATA[7]),
	.A1(Temp_Reg[7]),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[6]  (
	.SI(Temp_Reg[5]),
	.SE(n47),
	.RN(RST),
	.Q(Temp_Reg[6]),
	.D(n26),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[5]  (
	.SI(Temp_Reg[4]),
	.SE(n42),
	.RN(RST),
	.Q(Temp_Reg[5]),
	.D(n27),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[4]  (
	.SI(Temp_Reg[3]),
	.SE(n41),
	.RN(RST),
	.Q(Temp_Reg[4]),
	.D(n28),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[3]  (
	.SI(Temp_Reg[2]),
	.SE(n42),
	.RN(RST),
	.Q(Temp_Reg[3]),
	.D(n29),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[2]  (
	.SI(Temp_Reg[1]),
	.SE(n41),
	.RN(RST),
	.Q(Temp_Reg[2]),
	.D(n30),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[1]  (
	.SI(ser_data),
	.SE(n46),
	.RN(RST),
	.Q(Temp_Reg[1]),
	.D(n31),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[0]  (
	.SI(n35),
	.SE(n45),
	.RN(RST),
	.Q(ser_data),
	.D(n24),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Temp_Reg_reg[7]  (
	.SI(Temp_Reg[6]),
	.SE(n48),
	.RN(RST),
	.Q(Temp_Reg[7]),
	.D(n25),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \P_Counter_reg[2]  (
	.SI(P_Counter[1]),
	.SE(n47),
	.RN(RST),
	.QN(n35),
	.Q(P_Counter[2]),
	.D(n21),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \P_Counter_reg[0]  (
	.SI(test_si),
	.SE(n45),
	.RN(RST),
	.QN(n33),
	.Q(P_Counter[0]),
	.D(n23),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \P_Counter_reg[1]  (
	.SI(n33),
	.SE(n46),
	.RN(RST),
	.QN(n34),
	.Q(P_Counter[1]),
	.D(n22),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M ser_done_reg (
	.SI(Temp_Reg[7]),
	.SE(n48),
	.RN(RST),
	.QN(test_so),
	.Q(ser_done),
	.D(n20),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U35 (
	.Y(n39),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U36 (
	.Y(n40),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U37 (
	.Y(n41),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U38 (
	.Y(n42),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U39 (
	.Y(n43),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U40 (
	.Y(n44),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U41 (
	.Y(n45),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U42 (
	.Y(n46),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U43 (
	.Y(n47),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U44 (
	.Y(n48),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U45 (
	.Y(n49),
	.A(test_so), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_T_FSM_test_1 (
	Data_Valid, 
	PAR_EN, 
	ser_done, 
	CLK, 
	RST, 
	mux_sel, 
	Busy, 
	ser_en, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_O_RST3, 
	O_CLK3__L3_N2, 
	VDD, 
	VSS);
   input Data_Valid;
   input PAR_EN;
   input ser_done;
   input CLK;
   input RST;
   output [1:0] mux_sel;
   output Busy;
   output ser_en;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_O_RST3;
   input O_CLK3__L3_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire Busy_comb;
   wire n5;
   wire n6;
   wire n7;
   wire n2;
   wire n4;
   wire n8;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = n2 ;

   // Module instantiations
   INVX2M U4 (
	.Y(n2),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(ser_en),
	.B(current_state[2]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U6 (
	.Y(mux_sel[0]),
	.B(n2),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U8 (
	.Y(next_state[1]),
	.B0(mux_sel[1]),
	.A1N(n6),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U9 (
	.Y(next_state[0]),
	.B1(n7),
	.B0(current_state[1]),
	.A1(mux_sel[1]),
	.A0(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U10 (
	.Y(n7),
	.B0(ser_en),
	.A1(n2),
	.A0(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U11 (
	.Y(n6),
	.B(n8),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(mux_sel[1]),
	.A(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U13 (
	.Y(Busy_comb),
	.B0(mux_sel[1]),
	.A1(current_state[0]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n8),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(next_state[2]),
	.C(n5),
	.B(current_state[2]),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U16 (
	.Y(n5),
	.B0(n4),
	.A1N(PAR_EN),
	.A0(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(n15),
	.RN(FE_OFN4_O_RST3),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \current_state_reg[0]  (
	.SI(n12),
	.SE(n15),
	.RN(FE_OFN4_O_RST3),
	.QN(n4),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M Busy_reg (
	.SI(test_si),
	.SE(n14),
	.RN(RST),
	.QN(n12),
	.Q(Busy),
	.D(Busy_comb),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U17 (
	.Y(n13),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U18 (
	.Y(n14),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U19 (
	.Y(n15),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n8),
	.SE(n14),
	.RN(FE_OFN4_O_RST3),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_Parity_calc_test_1 (
	P_DATA, 
	Data_Valid, 
	PAR_TYPE, 
	PAR_EN, 
	CLK, 
	RST, 
	Busy, 
	par_bit, 
	test_si, 
	test_se, 
	FE_OFN4_O_RST3, 
	VDD, 
	VSS);
   input [7:0] P_DATA;
   input Data_Valid;
   input PAR_TYPE;
   input PAR_EN;
   input CLK;
   input RST;
   input Busy;
   output par_bit;
   input test_si;
   input test_se;
   input FE_OFN4_O_RST3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n19;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire [7:0] Data_draft;

   // Module instantiations
   NOR2BX2M U5 (
	.Y(n7),
	.B(Busy),
	.AN(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U6 (
	.Y(n9),
	.B1(n7),
	.B0(P_DATA[0]),
	.A1N(n7),
	.A0(Data_draft[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U7 (
	.Y(n10),
	.B1(n7),
	.B0(P_DATA[1]),
	.A1N(n7),
	.A0(Data_draft[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U8 (
	.Y(n11),
	.B1(n7),
	.B0(P_DATA[2]),
	.A1N(n7),
	.A0(Data_draft[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U9 (
	.Y(n12),
	.B1(n7),
	.B0(P_DATA[3]),
	.A1N(n7),
	.A0(Data_draft[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U10 (
	.Y(n13),
	.B1(n7),
	.B0(P_DATA[4]),
	.A1N(n7),
	.A0(Data_draft[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U11 (
	.Y(n14),
	.B1(n7),
	.B0(P_DATA[5]),
	.A1N(n7),
	.A0(Data_draft[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U12 (
	.Y(n15),
	.B1(n7),
	.B0(P_DATA[6]),
	.A1N(n7),
	.A0(Data_draft[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U13 (
	.Y(n16),
	.B1(n7),
	.B0(P_DATA[7]),
	.A1N(n7),
	.A0(Data_draft[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U14 (
	.Y(n5),
	.B(Data_draft[3]),
	.A(Data_draft[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U15 (
	.Y(n8),
	.B1(n19),
	.B0(n1),
	.A1N(n19),
	.A0N(par_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n19),
	.A(PAR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U17 (
	.Y(n1),
	.C(n4),
	.B(PAR_TYPE),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U18 (
	.Y(n4),
	.C(n5),
	.B(Data_draft[0]),
	.A(Data_draft[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U19 (
	.Y(n3),
	.C(n6),
	.B(Data_draft[4]),
	.A(Data_draft[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U20 (
	.Y(n6),
	.B(Data_draft[6]),
	.A(Data_draft[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M par_bit_reg (
	.SI(Data_draft[7]),
	.SE(n25),
	.RN(RST),
	.Q(par_bit),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[5]  (
	.SI(Data_draft[4]),
	.SE(n25),
	.RN(RST),
	.Q(Data_draft[5]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[1]  (
	.SI(Data_draft[0]),
	.SE(n27),
	.RN(RST),
	.Q(Data_draft[1]),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[4]  (
	.SI(Data_draft[3]),
	.SE(n24),
	.RN(FE_OFN4_O_RST3),
	.Q(Data_draft[4]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[0]  (
	.SI(test_si),
	.SE(n26),
	.RN(RST),
	.Q(Data_draft[0]),
	.D(n9),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[2]  (
	.SI(Data_draft[1]),
	.SE(n28),
	.RN(RST),
	.Q(Data_draft[2]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[7]  (
	.SI(Data_draft[6]),
	.SE(n24),
	.RN(FE_OFN4_O_RST3),
	.Q(Data_draft[7]),
	.D(n16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[3]  (
	.SI(Data_draft[2]),
	.SE(n23),
	.RN(RST),
	.Q(Data_draft[3]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Data_draft_reg[6]  (
	.SI(Data_draft[5]),
	.SE(n23),
	.RN(RST),
	.Q(Data_draft[6]),
	.D(n15),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U21 (
	.Y(n22),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U22 (
	.Y(n23),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U23 (
	.Y(n24),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U24 (
	.Y(n25),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U25 (
	.Y(n26),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U26 (
	.Y(n27),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U27 (
	.Y(n28),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_MUX_test_1 (
	mux_sel, 
	start_bit, 
	stop_bit, 
	ser_data, 
	par_bit, 
	CLK, 
	RST, 
	TX_OUT, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [1:0] mux_sel;
   input start_bit;
   input stop_bit;
   input ser_data;
   input par_bit;
   input CLK;
   input RST;
   output TX_OUT;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire out;
   wire n2;
   wire n3;
   wire n1;
   wire n5;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U4 (
	.Y(TX_OUT),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n5),
	.A(mux_sel[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U6 (
	.Y(out),
	.B1(n3),
	.B0(mux_sel[1]),
	.A1N(mux_sel[1]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U7 (
	.Y(n2),
	.B1(mux_sel[0]),
	.B0(LTIE_LTIELO_NET),
	.A1(n5),
	.A0(par_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U8 (
	.Y(n3),
	.B1(mux_sel[0]),
	.B0(ser_data),
	.A1(n5),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSX1M TX_OUT_reg (
	.SN(RST),
	.SI(test_si),
	.SE(test_se),
	.QN(n1),
	.D(out),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_RX_test_1 (
	CLK, 
	RST, 
	RX_IN, 
	parity_enable, 
	parity_type, 
	Prescale, 
	P_DATA, 
	data_valid, 
	parity_error, 
	framing_error, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN4_O_RST3, 
	O_CLK4__L3_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input RX_IN;
   input parity_enable;
   input parity_type;
   input [5:0] Prescale;
   output [7:0] P_DATA;
   output data_valid;
   output parity_error;
   output framing_error;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN4_O_RST3;
   input O_CLK4__L3_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire strt_glitch;
   wire strt_chk_en;
   wire edge_bit_en;
   wire deser_en;
   wire par_chk_en;
   wire stp_chk_en;
   wire dat_samp_en;
   wire sampled_bit;
   wire n5;
   wire n15;
   wire n26;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire [3:0] bit_count;
   wire [5:0] edge_count;

   // Module instantiations
   DLY1X1M U9 (
	.Y(n15),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U20 (
	.Y(n26),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U31 (
	.Y(n37),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U32 (
	.Y(n38),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U33 (
	.Y(n39),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U34 (
	.Y(n40),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U35 (
	.Y(n41),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U36 (
	.Y(n42),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U37 (
	.Y(n43),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   uart_rx_fsm_DATA_WIDTH8_test_1 U0_uart_fsm (
	.CLK(O_CLK4__L3_N1),
	.RST(FE_OFN4_O_RST3),
	.S_DATA(RX_IN),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		n26 }),
	.parity_enable(parity_enable),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.par_err(parity_error),
	.stp_err(framing_error),
	.strt_glitch(strt_glitch),
	.strt_chk_en(strt_chk_en),
	.edge_bit_en(edge_bit_en),
	.deser_en(deser_en),
	.par_chk_en(par_chk_en),
	.stp_chk_en(stp_chk_en),
	.dat_samp_en(dat_samp_en),
	.data_valid(data_valid),
	.test_so(test_so2),
	.test_se(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   edge_bit_counter_test_1 U0_edge_bit_counter (
	.CLK(CLK),
	.RST(FE_OFN4_O_RST3),
	.Enable(edge_bit_en),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.test_si2(test_si2),
	.test_si1(n5),
	.test_so1(test_so1),
	.test_se(n42),
	.O_CLK4__L3_N1(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   data_sampling_test_1 U0_data_sampling (
	.CLK(O_CLK4__L3_N1),
	.RST(FE_OFN4_O_RST3),
	.S_DATA(RX_IN),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		n26 }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.Enable(dat_samp_en),
	.sampled_bit(sampled_bit),
	.test_si(test_si1),
	.test_se(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_DATA_WIDTH8_test_1 U0_deserializer (
	.CLK(CLK),
	.RST(RST),
	.sampled_bit(sampled_bit),
	.Enable(deser_en),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.test_so(n5),
	.test_se(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   strt_chk_test_1 U0_strt_chk (
	.CLK(O_CLK4__L3_N1),
	.RST(FE_OFN4_O_RST3),
	.sampled_bit(sampled_bit),
	.Enable(strt_chk_en),
	.strt_glitch(strt_glitch),
	.test_si(framing_error),
	.test_se(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   par_chk_DATA_WIDTH8_test_1 U0_par_chk (
	.CLK(O_CLK4__L3_N1),
	.RST(FE_OFN4_O_RST3),
	.parity_type(parity_type),
	.sampled_bit(sampled_bit),
	.Enable(par_chk_en),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.par_err(parity_error),
	.test_si(edge_count[5]),
	.test_se(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   stp_chk_test_1 U0_stp_chk (
	.CLK(O_CLK4__L3_N1),
	.RST(FE_OFN4_O_RST3),
	.sampled_bit(sampled_bit),
	.Enable(stp_chk_en),
	.stp_err(framing_error),
	.test_si(parity_error),
	.test_se(n41), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module uart_rx_fsm_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	S_DATA, 
	Prescale, 
	parity_enable, 
	bit_count, 
	edge_count, 
	par_err, 
	stp_err, 
	strt_glitch, 
	strt_chk_en, 
	edge_bit_en, 
	deser_en, 
	par_chk_en, 
	stp_chk_en, 
	dat_samp_en, 
	data_valid, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input S_DATA;
   input [5:0] Prescale;
   input parity_enable;
   input [3:0] bit_count;
   input [5:0] edge_count;
   input par_err;
   input stp_err;
   input strt_glitch;
   output strt_chk_en;
   output edge_bit_en;
   output deser_en;
   output par_chk_en;
   output stp_chk_en;
   output dat_samp_en;
   output data_valid;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \sub_41/carry[5] ;
   wire \sub_41/carry[4] ;
   wire \sub_41/carry[3] ;
   wire n2;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n58;
   wire n59;
   wire n69;
   wire n71;
   wire [5:0] check_edge;
   wire [5:0] error_check_edge;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign error_check_edge[0] = Prescale[0] ;
   assign test_so = n33 ;

   // Module instantiations
   OR2X2M U5 (
	.Y(n5),
	.B(n54),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n17),
	.B(n2),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(n6),
	.B(Prescale[2]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U8 (
	.Y(dat_samp_en),
	.B(n10),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U9 (
	.Y(stp_chk_en),
	.B(n11),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U10 (
	.Y(strt_chk_en),
	.B(n10),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U11 (
	.Y(n10),
	.B0(n33),
	.A1(n40),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U13 (
	.Y(n23),
	.B1(n14),
	.B0(deser_en),
	.A1N(S_DATA),
	.A0N(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n25),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U15 (
	.Y(edge_bit_en),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U16 (
	.Y(n11),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n39),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U18 (
	.Y(n29),
	.C(n32),
	.B(n31),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BXLM U19 (
	.Y(n30),
	.C(stp_chk_en),
	.B(bit_count[3]),
	.AN(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U20 (
	.Y(deser_en),
	.C(current_state[2]),
	.B(n39),
	.AN(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n33),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BXLM U22 (
	.Y(next_state[2]),
	.C(n13),
	.B(n12),
	.AN(stp_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BXLM U23 (
	.Y(n13),
	.C(n15),
	.B(deser_en),
	.AN(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U24 (
	.Y(n16),
	.D(n45),
	.C(n44),
	.B(n43),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U25 (
	.Y(n19),
	.C(bit_count[3]),
	.B(strt_glitch),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1XLM U26 (
	.Y(check_edge[1]),
	.B0(n5),
	.A1N(Prescale[1]),
	.A0N(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U27 (
	.Y(n38),
	.B(n25),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U28 (
	.Y(n28),
	.C(n36),
	.B(n35),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U29 (
	.Y(n24),
	.C(n2),
	.B(current_state[1]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n9),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U32 (
	.Y(error_check_edge[1]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U33 (
	.Y(error_check_edge[5]),
	.B(\sub_41/carry[5] ),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U34 (
	.Y(\sub_41/carry[5] ),
	.B(\sub_41/carry[4] ),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U35 (
	.Y(error_check_edge[4]),
	.B(Prescale[4]),
	.A(\sub_41/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U36 (
	.Y(\sub_41/carry[4] ),
	.B(\sub_41/carry[3] ),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U37 (
	.Y(error_check_edge[3]),
	.B(n52),
	.A(\sub_41/carry[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U38 (
	.Y(\sub_41/carry[3] ),
	.B(Prescale[1]),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U39 (
	.Y(error_check_edge[2]),
	.B(Prescale[2]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U41 (
	.Y(check_edge[2]),
	.B0(n6),
	.A1(Prescale[2]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U42 (
	.Y(n7),
	.B(n9),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U43 (
	.Y(check_edge[3]),
	.B0(n7),
	.A1(n9),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U44 (
	.Y(check_edge[4]),
	.B(n7),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(check_edge[5]),
	.B(n71),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U47 (
	.Y(par_chk_en),
	.B(n11),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U48 (
	.Y(n15),
	.A(parity_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U49 (
	.Y(n12),
	.D(n17),
	.C(n16),
	.B(bit_count[0]),
	.A(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U50 (
	.Y(next_state[1]),
	.B0(n11),
	.A1(n18),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U51 (
	.Y(n18),
	.B0(current_state[1]),
	.A2(n19),
	.A1(n16),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U52 (
	.Y(next_state[0]),
	.C0(n23),
	.B0(n22),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U53 (
	.Y(n14),
	.C(bit_count[3]),
	.B(n25),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U54 (
	.Y(n22),
	.D(n29),
	.C(n28),
	.B(n27),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U55 (
	.Y(n32),
	.B(edge_count[5]),
	.A(error_check_edge[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n31),
	.B(edge_count[4]),
	.A(error_check_edge[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n36),
	.B(edge_count[1]),
	.A(error_check_edge[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(n35),
	.B(edge_count[0]),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n34),
	.B(error_check_edge[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U60 (
	.Y(n27),
	.B(error_check_edge[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U61 (
	.Y(n26),
	.S0(n53),
	.B(n38),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U62 (
	.Y(n37),
	.B(n25),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U63 (
	.Y(n21),
	.B(n33),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U64 (
	.Y(n20),
	.S0(n2),
	.B(n41),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U65 (
	.Y(n41),
	.D(n25),
	.C(n16),
	.B(strt_glitch),
	.AN(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U66 (
	.Y(n45),
	.D(n49),
	.C(n48),
	.B(n47),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U67 (
	.Y(n49),
	.B(check_edge[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U68 (
	.Y(n48),
	.B(check_edge[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U69 (
	.Y(n47),
	.B(check_edge[5]),
	.A(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U70 (
	.Y(n46),
	.B(check_edge[1]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(n44),
	.B(bit_count[1]),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U72 (
	.Y(n43),
	.B(check_edge[4]),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U73 (
	.Y(n42),
	.B(n69),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U74 (
	.Y(data_valid),
	.C(par_err),
	.B(stp_err),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U75 (
	.Y(n40),
	.A(S_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n39),
	.SE(n58),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n2),
	.SE(n59),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U40 (
	.Y(n52),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U45 (
	.Y(n53),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U76 (
	.Y(n54),
	.A(error_check_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U77 (
	.Y(n55),
	.A(error_check_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U80 (
	.Y(n58),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U81 (
	.Y(n59),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U92 (
	.Y(n69),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U94 (
	.Y(n8),
	.B(n7),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U95 (
	.Y(n71),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \current_state_reg[0]  (
	.SI(strt_glitch),
	.SE(n58),
	.RN(RST),
	.Q(n2),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module edge_bit_counter_test_1 (
	CLK, 
	RST, 
	Enable, 
	Prescale, 
	bit_count, 
	edge_count, 
	test_si2, 
	test_si1, 
	test_so1, 
	test_se, 
	O_CLK4__L3_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input Enable;
   input [5:0] Prescale;
   output [3:0] bit_count;
   output [5:0] edge_count;
   input test_si2;
   input test_si1;
   output test_so1;
   input test_se;
   input O_CLK4__L3_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire n53;
   wire n54;
   wire n56;
   wire n57;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire n4;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire \add_31/carry[5] ;
   wire \add_31/carry[4] ;
   wire \add_31/carry[3] ;
   wire \add_31/carry[2] ;
   wire n1;
   wire n52;
   wire n6;
   wire n55;
   wire n22;
   wire n24;
   wire n26;
   wire n58;
   wire n30;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n62;
   wire n63;
   wire n64;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n75;
   wire n76;
   wire n7;
   wire n21;
   wire n25;
   wire n28;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U3 (
	.Y(edge_count[5]),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(N25),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U9 (
	.Y(n6),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U10 (
	.Y(edge_count[4]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X1M U11 (
	.Y(n10),
	.B(n76),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U14 (
	.Y(n22),
	.A(test_so1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U15 (
	.Y(edge_count[2]),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U16 (
	.Y(n24),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U17 (
	.Y(n26),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U18 (
	.Y(edge_count[1]),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(n34),
	.B(Prescale[2]),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U22 (
	.Y(n33),
	.B(N25),
	.AN(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U23 (
	.Y(N31),
	.D(n43),
	.C(n44),
	.B(n45),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U24 (
	.Y(n39),
	.B(edge_count[0]),
	.AN(N25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U25 (
	.Y(n38),
	.B(N25),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U26 (
	.Y(n14),
	.C(Enable),
	.B(n47),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U29 (
	.Y(n47),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U30 (
	.Y(n50),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(n13),
	.B(N31),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U32 (
	.Y(n16),
	.B0(n13),
	.A1(Enable),
	.A0(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U33 (
	.Y(N20),
	.B(n47),
	.AN(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U34 (
	.Y(N21),
	.B(n47),
	.AN(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U35 (
	.Y(N22),
	.B(n47),
	.AN(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U36 (
	.Y(N23),
	.B(n47),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U37 (
	.Y(n20),
	.B1(n47),
	.B0(n48),
	.A2(n13),
	.A1(n76),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U38 (
	.Y(n18),
	.B1(n1),
	.B0(n15),
	.A2(n49),
	.A1(bit_count[2]),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U39 (
	.Y(n15),
	.B0N(n16),
	.A1(n49),
	.A0(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U40 (
	.Y(n19),
	.B1(n14),
	.B0(bit_count[1]),
	.A1(n49),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U41 (
	.Y(N24),
	.B(n47),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U42 (
	.Y(n30),
	.B(edge_count[5]),
	.A(\add_31/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U43 (
	.Y(N19),
	.B(n47),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U44 (
	.Y(n17),
	.B1(n4),
	.B0(n11),
	.A2(n50),
	.A1(n10),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3XLM U45 (
	.Y(n9),
	.C(n4),
	.B(bit_count[2]),
	.A(N31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U46 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U47 (
	.Y(n12),
	.B0(n50),
	.A1N(n1),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U48 (
	.S(N8),
	.CO(\add_31/carry[2] ),
	.B(edge_count[0]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U49 (
	.S(N9),
	.CO(\add_31/carry[3] ),
	.B(\add_31/carry[2] ),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U50 (
	.S(N10),
	.CO(\add_31/carry[4] ),
	.B(\add_31/carry[3] ),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U51 (
	.S(N11),
	.CO(\add_31/carry[5] ),
	.B(\add_31/carry[4] ),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n49),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U54 (
	.Y(n37),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U55 (
	.Y(N26),
	.B0(n33),
	.A1N(Prescale[1]),
	.A0N(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U56 (
	.Y(N27),
	.B0(n34),
	.A1(Prescale[2]),
	.A0(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U57 (
	.Y(n35),
	.B(n37),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U58 (
	.Y(N28),
	.B0(n35),
	.A1(n37),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U59 (
	.Y(N29),
	.B(n35),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U61 (
	.Y(N30),
	.B(n75),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U62 (
	.Y(n42),
	.B1(n38),
	.B0(edge_count[1]),
	.A1N(N26),
	.A0(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U63 (
	.Y(n41),
	.B1(n39),
	.B0(N26),
	.A1N(edge_count[1]),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U64 (
	.Y(n40),
	.B(edge_count[5]),
	.A(N30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U65 (
	.Y(n46),
	.C(n40),
	.B(n41),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U66 (
	.Y(n45),
	.B(edge_count[4]),
	.A(N29), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U67 (
	.Y(n44),
	.B(edge_count[2]),
	.A(N27), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U68 (
	.Y(n43),
	.B(edge_count[3]),
	.A(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \bit_count_reg[3]  (
	.SI(bit_count[2]),
	.SE(n68),
	.RN(RST),
	.QN(n4),
	.Q(bit_count[3]),
	.D(n17),
	.CK(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[1]  (
	.SI(edge_count[0]),
	.SE(n64),
	.RN(RST),
	.Q(n57),
	.D(N20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[5]  (
	.SI(edge_count[4]),
	.SE(n71),
	.RN(RST),
	.Q(n53),
	.D(N24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[4]  (
	.SI(edge_count[3]),
	.SE(n70),
	.RN(RST),
	.Q(n54),
	.D(N23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U60 (
	.Y(n62),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U69 (
	.Y(n63),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U70 (
	.Y(n64),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U72 (
	.Y(n66),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U73 (
	.Y(n67),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U74 (
	.Y(n68),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U75 (
	.Y(n69),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U76 (
	.Y(n70),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U77 (
	.Y(n71),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U82 (
	.Y(n36),
	.B(n35),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U83 (
	.Y(n75),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U84 (
	.Y(n76),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \edge_count_reg[3]  (
	.SI(test_si2),
	.SE(n69),
	.RN(RST),
	.Q(n55),
	.D(N22),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \edge_count_reg[0]  (
	.SI(n4),
	.SE(n71),
	.RN(RST),
	.Q(n58),
	.D(N19),
	.CK(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \bit_count_reg[1]  (
	.SI(n48),
	.SE(n63),
	.RN(RST),
	.Q(n52),
	.D(n19),
	.CK(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \bit_count_reg[2]  (
	.SI(n49),
	.SE(n70),
	.RN(RST),
	.QN(n1),
	.D(n18),
	.CK(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX2M \bit_count_reg[0]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(test_si1),
	.SE(n64),
	.RN(RST),
	.QN(n48),
	.Q(bit_count[0]),
	.D(n20),
	.CK(O_CLK4__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \edge_count_reg[2]  (
	.SI(edge_count[1]),
	.SE(n63),
	.RN(RST),
	.Q(n56),
	.D(N21),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U7 (
	.Y(bit_count[2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U12 (
	.Y(n7),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U13 (
	.Y(bit_count[1]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U19 (
	.Y(n21),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX8M U20 (
	.Y(test_so1),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U53 (
	.Y(n25),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U94 (
	.Y(edge_count[3]),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U95 (
	.Y(n28),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U96 (
	.Y(edge_count[0]),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampling_test_1 (
	CLK, 
	RST, 
	S_DATA, 
	Prescale, 
	edge_count, 
	Enable, 
	sampled_bit, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input S_DATA;
   input [5:0] Prescale;
   input [5:0] edge_count;
   input Enable;
   output sampled_bit;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N58;
   wire n19;
   wire n20;
   wire n21;
   wire \add_21/carry[4] ;
   wire \add_21/carry[3] ;
   wire \add_21/carry[2] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n40;
   wire n41;
   wire n44;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n53;
   wire [4:0] half_edges;
   wire [4:0] half_edges_p1;
   wire [4:0] half_edges_n1;
   wire [2:0] Samples;

   // Module instantiations
   INVX2M U3 (
	.Y(half_edges[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U4 (
	.Y(n17),
	.D(n37),
	.C(n36),
	.B(n35),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U5 (
	.Y(n12),
	.D(n16),
	.C(n15),
	.B(n14),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n6),
	.B(half_edges[0]),
	.A(half_edges[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U7 (
	.Y(half_edges[1]),
	.B0(n49),
	.A1(Prescale[2]),
	.A0(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U8 (
	.Y(half_edges[2]),
	.B0(n3),
	.A1(n5),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(half_edges[3]),
	.B(n3),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U11 (
	.Y(n3),
	.B(n5),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U12 (
	.Y(n33),
	.B(Enable),
	.A(Samples[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U13 (
	.Y(n26),
	.B(Enable),
	.A(Samples[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U14 (
	.Y(n32),
	.B(edge_count[1]),
	.A(half_edges[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U15 (
	.Y(n31),
	.B(edge_count[0]),
	.A(half_edges[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U16 (
	.Y(n10),
	.B(Enable),
	.A(Samples[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U17 (
	.Y(n37),
	.C(n16),
	.B(edge_count[5]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U19 (
	.Y(n9),
	.A(half_edges[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U20 (
	.S(half_edges_p1[2]),
	.CO(\add_21/carry[3] ),
	.B(\add_21/carry[2] ),
	.A(half_edges[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U21 (
	.S(half_edges_p1[3]),
	.CO(\add_21/carry[4] ),
	.B(\add_21/carry[3] ),
	.A(half_edges[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U22 (
	.S(half_edges_p1[1]),
	.CO(\add_21/carry[2] ),
	.B(half_edges[0]),
	.A(half_edges[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n5),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U25 (
	.Y(half_edges[4]),
	.B(n53),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U26 (
	.Y(half_edges_p1[4]),
	.B(half_edges[4]),
	.A(\add_21/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U27 (
	.Y(half_edges_n1[1]),
	.B0(n6),
	.A1(half_edges[1]),
	.A0(half_edges[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U28 (
	.Y(n7),
	.B(n9),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U29 (
	.Y(half_edges_n1[2]),
	.B0(n7),
	.A1(n9),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U30 (
	.Y(half_edges_n1[3]),
	.B(n7),
	.A(half_edges[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U31 (
	.Y(n8),
	.B(n7),
	.A(half_edges[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(half_edges_n1[4]),
	.B(n8),
	.A(half_edges[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U33 (
	.Y(n21),
	.S0(n12),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U34 (
	.Y(n16),
	.B(edge_count[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U35 (
	.Y(n14),
	.B(n17),
	.A(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U36 (
	.Y(n13),
	.D(n24),
	.C(n23),
	.B(n22),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U37 (
	.Y(n24),
	.B(half_edges_p1[1]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U38 (
	.Y(n23),
	.B(half_edges_p1[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U39 (
	.Y(n22),
	.B(half_edges_p1[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n18),
	.B(half_edges_p1[4]),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U41 (
	.Y(n20),
	.S0(n15),
	.B(n11),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U42 (
	.Y(n15),
	.D(n30),
	.C(n29),
	.B(n28),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U43 (
	.Y(n30),
	.D(n32),
	.C(n31),
	.B(n17),
	.A(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U44 (
	.Y(n29),
	.B(half_edges[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U45 (
	.Y(n28),
	.B(half_edges[4]),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U46 (
	.Y(n25),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U47 (
	.Y(n27),
	.B(half_edges[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U48 (
	.Y(n19),
	.S0(n17),
	.B(n11),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n38),
	.B(edge_count[4]),
	.A(half_edges_n1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U51 (
	.Y(n36),
	.B(half_edges_n1[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U52 (
	.Y(n35),
	.B(half_edges_n1[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U53 (
	.Y(n34),
	.B(half_edges_n1[1]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U54 (
	.Y(n11),
	.B(Enable),
	.A(S_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX1M U55 (
	.Y(N58),
	.B0N(Enable),
	.A1(n41),
	.A0(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U9 (
	.Y(n44),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U58 (
	.Y(n46),
	.B(Prescale[1]),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U59 (
	.Y(n47),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U60 (
	.Y(n48),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U61 (
	.Y(n49),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U65 (
	.Y(n4),
	.B(n3),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U66 (
	.Y(n53),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M sampled_bit_reg (
	.SI(Samples[2]),
	.SE(n48),
	.RN(RST),
	.Q(sampled_bit),
	.D(N58),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Samples_reg[2]  (
	.SI(Samples[1]),
	.SE(n47),
	.RN(RST),
	.Q(Samples[2]),
	.D(n21),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX2M \Samples_reg[0]  (
	.SI(test_si),
	.SE(n47),
	.RN(RST),
	.Q(Samples[0]),
	.D(n19),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX2M \Samples_reg[1]  (
	.SI(Samples[0]),
	.SE(n48),
	.RN(RST),
	.Q(Samples[1]),
	.D(n20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U56 (
	.Y(n41),
	.B0(Samples[2]),
	.A1(Samples[1]),
	.A0(Samples[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U73 (
	.Y(n40),
	.B(Samples[1]),
	.A(Samples[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	sampled_bit, 
	Enable, 
	edge_count, 
	Prescale, 
	P_DATA, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input sampled_bit;
   input Enable;
   input [5:0] edge_count;
   input [5:0] Prescale;
   output [7:0] P_DATA;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N1;
   wire N2;
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire n1;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n44;

   assign test_so = n27 ;

   // Module instantiations
   INVX2M U3 (
	.Y(N1),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U4 (
	.Y(n6),
	.B(Prescale[2]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U5 (
	.Y(n5),
	.B(N1),
	.AN(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U6 (
	.Y(n18),
	.B(N1),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U7 (
	.Y(n19),
	.B(edge_count[0]),
	.AN(N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U10 (
	.Y(n34),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U11 (
	.Y(n11),
	.B1(n32),
	.B0(n1),
	.A1(n33),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U12 (
	.Y(n12),
	.B1(n31),
	.B0(n1),
	.A1(n32),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U13 (
	.Y(n13),
	.B1(n30),
	.B0(n1),
	.A1(n31),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U14 (
	.Y(n14),
	.B1(n29),
	.B0(n1),
	.A1(n30),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U15 (
	.Y(n15),
	.B1(n28),
	.B0(n1),
	.A1(n29),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U16 (
	.Y(n16),
	.B1(n27),
	.B0(n1),
	.A1(n28),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U17 (
	.Y(n17),
	.B1(n27),
	.B0(n34),
	.A1N(n34),
	.A0N(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U18 (
	.Y(n10),
	.B1(n33),
	.B0(n1),
	.A1N(n1),
	.A0N(P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U20 (
	.Y(n1),
	.B(Enable),
	.A(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n32),
	.A(P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n28),
	.A(P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n27),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n31),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n33),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n30),
	.A(P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n29),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n9),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U29 (
	.Y(N2),
	.B0(n5),
	.A1N(Prescale[1]),
	.A0N(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U30 (
	.Y(N3),
	.B0(n6),
	.A1(Prescale[2]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U31 (
	.Y(n7),
	.B(n9),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U32 (
	.Y(N4),
	.B0(n7),
	.A1(n9),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U33 (
	.Y(N5),
	.B(n7),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U35 (
	.Y(N6),
	.B(n44),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U36 (
	.Y(n22),
	.B1(n18),
	.B0(edge_count[1]),
	.A1N(N2),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U37 (
	.Y(n21),
	.B1(n19),
	.B0(N2),
	.A1N(edge_count[1]),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U38 (
	.Y(n20),
	.B(edge_count[5]),
	.A(N6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U39 (
	.Y(n26),
	.C(n20),
	.B(n21),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n25),
	.B(edge_count[4]),
	.A(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(n24),
	.B(edge_count[2]),
	.A(N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n23),
	.B(edge_count[3]),
	.A(N4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U43 (
	.Y(N7),
	.D(n23),
	.C(n24),
	.B(n25),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[0]  (
	.SI(sampled_bit),
	.SE(n39),
	.RN(RST),
	.Q(P_DATA[0]),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[5]  (
	.SI(n30),
	.SE(n41),
	.RN(RST),
	.Q(P_DATA[5]),
	.D(n15),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[1]  (
	.SI(P_DATA[0]),
	.SE(n40),
	.RN(RST),
	.Q(P_DATA[1]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[4]  (
	.SI(n31),
	.SE(n38),
	.RN(RST),
	.Q(P_DATA[4]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[7]  (
	.SI(n28),
	.SE(n38),
	.RN(RST),
	.Q(P_DATA[7]),
	.D(n17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[3]  (
	.SI(n32),
	.SE(n37),
	.RN(RST),
	.Q(P_DATA[3]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[6]  (
	.SI(n29),
	.SE(n37),
	.RN(RST),
	.Q(P_DATA[6]),
	.D(n16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[2]  (
	.SI(n33),
	.SE(n41),
	.RN(RST),
	.Q(P_DATA[2]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U34 (
	.Y(n36),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U44 (
	.Y(n37),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U45 (
	.Y(n38),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U46 (
	.Y(n39),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U47 (
	.Y(n40),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U48 (
	.Y(n41),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U51 (
	.Y(n8),
	.B(n7),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U52 (
	.Y(n44),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module strt_chk_test_1 (
	CLK, 
	RST, 
	sampled_bit, 
	Enable, 
	strt_glitch, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input sampled_bit;
   input Enable;
   output strt_glitch;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;

   // Module instantiations
   AO2B2XLM U2 (
	.Y(n1),
	.B1(Enable),
	.B0(sampled_bit),
	.A1N(Enable),
	.A0(strt_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M strt_glitch_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(strt_glitch),
	.D(n1),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module par_chk_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	parity_type, 
	sampled_bit, 
	Enable, 
	P_DATA, 
	par_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input parity_type;
   input sampled_bit;
   input Enable;
   input [7:0] P_DATA;
   output par_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n10;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;

   // Module instantiations
   BUFX10M U2 (
	.Y(par_err),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U3 (
	.Y(n8),
	.B1(n9),
	.B0(n1),
	.A1N(n9),
	.A0N(par_err), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U4 (
	.Y(n1),
	.C(n5),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n9),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(n5),
	.B(parity_type),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U7 (
	.Y(n4),
	.C(n6),
	.B(P_DATA[4]),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U8 (
	.Y(n6),
	.B(P_DATA[6]),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U9 (
	.Y(n3),
	.C(n7),
	.B(P_DATA[0]),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n7),
	.B(P_DATA[2]),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M par_err_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(n10),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stp_chk_test_1 (
	CLK, 
	RST, 
	sampled_bit, 
	Enable, 
	stp_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input sampled_bit;
   input Enable;
   output stp_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n4;
   wire n2;
   wire n3;

   // Module instantiations
   BUFX10M U2 (
	.Y(stp_err),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U3 (
	.Y(n2),
	.B1(n3),
	.B0(sampled_bit),
	.A1N(n3),
	.A0N(stp_err), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U4 (
	.Y(n3),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M stp_err_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(n4),
	.D(n2),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYSTEM_CTRL_BYTE8_test_1 (
	ALU_OUT, 
	ALU_OUT_VLD, 
	RX_P_DATA, 
	RX_D_VLD, 
	FIFO_FULL, 
	RdData, 
	RdData_Valid, 
	CLK, 
	RST, 
	ALU_EN, 
	ALU_FUN, 
	CLK_EN, 
	Address, 
	WrEn, 
	RdEn, 
	WrData, 
	TX_P_Data, 
	TX_D_VLD, 
	clk_div_en, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN3_O_RST2, 
	O_CLK1__L5_N7, 
	VDD, 
	VSS);
   input [15:0] ALU_OUT;
   input ALU_OUT_VLD;
   input [7:0] RX_P_DATA;
   input RX_D_VLD;
   input FIFO_FULL;
   input [7:0] RdData;
   input RdData_Valid;
   input CLK;
   input RST;
   output ALU_EN;
   output [3:0] ALU_FUN;
   output CLK_EN;
   output [3:0] Address;
   output WrEn;
   output RdEn;
   output [7:0] WrData;
   output [7:0] TX_P_Data;
   output TX_D_VLD;
   output clk_div_en;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN3_O_RST2;
   input O_CLK1__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire n99;
   wire n100;
   wire frame_flag;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n105;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire [3:0] current_state;
   wire [3:0] next_state;
   wire [3:0] Address_seq;

   assign test_so = n6 ;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U16 (
	.Y(n41),
	.B0(n34),
	.A2(n47),
	.A1(n92),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U53 (
	.Y(n53),
	.C(n50),
	.B(n6),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(ALU_FUN[3]),
	.B(n20),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(ALU_FUN[1]),
	.B(n20),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(ALU_FUN[0]),
	.B(n20),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U8 (
	.Y(n72),
	.B(RX_D_VLD),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U9 (
	.Y(n46),
	.C(RX_P_DATA[0]),
	.B(n91),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n3),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U12 (
	.Y(n51),
	.B0(n55),
	.A1(n88),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n6),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n5),
	.A(frame_flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U15 (
	.Y(n47),
	.B(RX_P_DATA[4]),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U19 (
	.Y(Address[3]),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U20 (
	.Y(n99),
	.B1(n72),
	.B0(n94),
	.A1N(Address_seq[3]),
	.A0(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U21 (
	.Y(Address[2]),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U22 (
	.Y(n100),
	.B1(n72),
	.B0(n95),
	.A1N(Address_seq[2]),
	.A0(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(ALU_FUN[2]),
	.B(n20),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(WrEn),
	.B(n52),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U25 (
	.Y(n40),
	.B(n37),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U26 (
	.Y(n30),
	.B(current_state[1]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U27 (
	.Y(n98),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n97),
	.A(RX_P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n91),
	.A(RX_P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n92),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U31 (
	.Y(n20),
	.A(ALU_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U32 (
	.Y(n52),
	.B(n22),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U33 (
	.Y(n21),
	.A(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U34 (
	.Y(ALU_EN),
	.B(n68),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U35 (
	.Y(n68),
	.B(n30),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U36 (
	.Y(n71),
	.B0(n73),
	.A1(n22),
	.A0(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U37 (
	.Y(n73),
	.D(n76),
	.C(n70),
	.B(n67),
	.AN(CLK_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U38 (
	.Y(n76),
	.B0(n78),
	.A1(n98),
	.A0(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U39 (
	.Y(n77),
	.B(n37),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U40 (
	.Y(n67),
	.C(n79),
	.B(n70),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U41 (
	.Y(n79),
	.C(n86),
	.B(CLK_EN),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U42 (
	.Y(CLK_EN),
	.B(n50),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U43 (
	.Y(n39),
	.B(n29),
	.AN(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n22),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n86),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U46 (
	.Y(n45),
	.B(n30),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U47 (
	.Y(n55),
	.B(n70),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n18),
	.A(FIFO_FULL), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U49 (
	.Y(n56),
	.B(n50),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U50 (
	.Y(WrData[0]),
	.B(n21),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U51 (
	.Y(WrData[1]),
	.B(n21),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U52 (
	.Y(WrData[2]),
	.B(n21),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U54 (
	.Y(WrData[3]),
	.B(n21),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U55 (
	.Y(WrData[4]),
	.B(n21),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U56 (
	.Y(WrData[5]),
	.B(n21),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U57 (
	.Y(WrData[6]),
	.B(n21),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U58 (
	.Y(n88),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U59 (
	.Y(n17),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U60 (
	.Y(n28),
	.B(n24),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U61 (
	.Y(RdEn),
	.B(n98),
	.AN(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U62 (
	.Y(next_state[1]),
	.C0(n38),
	.B1(n37),
	.B0(n98),
	.A1(n36),
	.A0(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U63 (
	.Y(n90),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U64 (
	.Y(n38),
	.C0(n40),
	.B0(n28),
	.A1(n98),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U65 (
	.Y(next_state[3]),
	.B0(n20),
	.A1N(n88),
	.A0N(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U66 (
	.Y(n24),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U67 (
	.Y(n49),
	.C(n95),
	.B(n91),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U68 (
	.Y(n87),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U69 (
	.Y(n23),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U72 (
	.Y(n35),
	.B(current_state[3]),
	.AN(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U73 (
	.Y(n50),
	.C(current_state[3]),
	.B(n30),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U74 (
	.Y(n80),
	.B(current_state[3]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U75 (
	.Y(n70),
	.C(current_state[1]),
	.B(n3),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U76 (
	.Y(n96),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U77 (
	.Y(n29),
	.C(current_state[1]),
	.B(n35),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U78 (
	.Y(n95),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U79 (
	.Y(n74),
	.C(n4),
	.B(n89),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U80 (
	.Y(n78),
	.C(current_state[1]),
	.B(n3),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U81 (
	.Y(n89),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U82 (
	.Y(n94),
	.A(RX_P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U84 (
	.Y(n37),
	.B(n4),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U86 (
	.Y(Address[0]),
	.C0(n75),
	.B1(n74),
	.B0(n98),
	.A1(n72),
	.A0(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U87 (
	.Y(n75),
	.B0(Address_seq[0]),
	.A1(n73),
	.A0(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U89 (
	.Y(Address[1]),
	.B1(n72),
	.B0(n96),
	.A1N(Address_seq[1]),
	.A0(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U90 (
	.Y(n69),
	.B(n18),
	.A(RdData_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U91 (
	.Y(n81),
	.B0(Address[3]),
	.A1(Address_seq[3]),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U92 (
	.Y(n82),
	.B0(Address[2]),
	.A1(Address_seq[2]),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U93 (
	.Y(n66),
	.C0(n63),
	.B1(n6),
	.B0(ALU_OUT[8]),
	.A1(n5),
	.A0(ALU_OUT[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U94 (
	.Y(TX_P_Data[0]),
	.C(n52),
	.B(n65),
	.AN(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U95 (
	.Y(n64),
	.D(n68),
	.C(n37),
	.B(n67),
	.AN(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U96 (
	.Y(n65),
	.B1(n24),
	.B0(RdData[0]),
	.A1N(n50),
	.A0N(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U97 (
	.Y(TX_P_Data[1]),
	.B0(n62),
	.A1N(n53),
	.A0N(ALU_OUT[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U98 (
	.Y(n62),
	.B1(n56),
	.B0(ALU_OUT[9]),
	.A1(n55),
	.A0(RdData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U99 (
	.Y(TX_P_Data[2]),
	.B0(n61),
	.A1N(n53),
	.A0N(ALU_OUT[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U100 (
	.Y(n61),
	.B1(n56),
	.B0(ALU_OUT[10]),
	.A1(n55),
	.A0(RdData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U101 (
	.Y(TX_P_Data[3]),
	.B0(n60),
	.A1N(n53),
	.A0N(ALU_OUT[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U102 (
	.Y(n60),
	.B1(n56),
	.B0(ALU_OUT[11]),
	.A1(n55),
	.A0(RdData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U103 (
	.Y(TX_P_Data[4]),
	.B0(n59),
	.A1N(n53),
	.A0N(ALU_OUT[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U104 (
	.Y(n59),
	.B1(n56),
	.B0(ALU_OUT[12]),
	.A1(n55),
	.A0(RdData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U105 (
	.Y(TX_P_Data[5]),
	.B0(n58),
	.A1N(n53),
	.A0N(ALU_OUT[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U106 (
	.Y(n58),
	.B1(n56),
	.B0(ALU_OUT[13]),
	.A1(n55),
	.A0(RdData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U107 (
	.Y(TX_P_Data[6]),
	.B0(n57),
	.A1N(n53),
	.A0N(ALU_OUT[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U108 (
	.Y(n57),
	.B1(n56),
	.B0(ALU_OUT[14]),
	.A1(n55),
	.A0(RdData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U109 (
	.Y(TX_P_Data[7]),
	.B0(n54),
	.A1N(n53),
	.A0N(ALU_OUT[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U110 (
	.Y(n54),
	.B1(n56),
	.B0(ALU_OUT[15]),
	.A1(n55),
	.A0(RdData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U111 (
	.Y(WrData[7]),
	.B(n21),
	.AN(RX_P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U112 (
	.Y(n25),
	.B(n17),
	.A(frame_flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U113 (
	.Y(n63),
	.B(n18),
	.A(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U114 (
	.Y(n84),
	.B1(Address_seq[0]),
	.B0(n37),
	.A1(n86),
	.A0(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U115 (
	.Y(n83),
	.B0(Address[1]),
	.A1(Address_seq[1]),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U116 (
	.Y(n85),
	.B1(n5),
	.B0(TX_D_VLD),
	.A2(n51),
	.A1(n6),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U117 (
	.Y(TX_D_VLD),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U118 (
	.Y(next_state[2]),
	.C0(n27),
	.B0(n26),
	.A1(n19),
	.A0(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U119 (
	.Y(n19),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U120 (
	.Y(n27),
	.C(n28),
	.B(RdEn),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U121 (
	.Y(n26),
	.B1(n31),
	.B0(n87),
	.A2(current_state[2]),
	.A1(n25),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U122 (
	.Y(n31),
	.B0(n34),
	.A2(n33),
	.A1(n91),
	.A0(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U123 (
	.Y(n33),
	.B(RX_P_DATA[2]),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U124 (
	.Y(n32),
	.C(RX_P_DATA[0]),
	.B(n92),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U125 (
	.Y(n34),
	.D(n48),
	.C(RX_P_DATA[6]),
	.B(n97),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U126 (
	.Y(n48),
	.C(n105),
	.B(RX_P_DATA[5]),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U127 (
	.Y(n36),
	.D(RX_D_VLD),
	.C(n45),
	.B(RX_P_DATA[3]),
	.A(RX_P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U128 (
	.Y(n93),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U129 (
	.Y(next_state[0]),
	.C(n43),
	.B(n29),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X2M U130 (
	.Y(n43),
	.C(n3),
	.B(RX_D_VLD),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U131 (
	.Y(n42),
	.B0(n87),
	.A1(n41),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U132 (
	.Y(n44),
	.D(n96),
	.C(RX_P_DATA[0]),
	.B(n92),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n89),
	.SE(n108),
	.RN(FE_OFN3_O_RST2),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[3]  (
	.SI(current_state[2]),
	.SE(n109),
	.RN(FE_OFN3_O_RST2),
	.Q(current_state[3]),
	.D(next_state[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(Address_seq[3]),
	.SE(n109),
	.RN(FE_OFN3_O_RST2),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n4),
	.SE(n110),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M frame_flag_reg (
	.SI(current_state[3]),
	.SE(n110),
	.RN(FE_OFN3_O_RST2),
	.Q(frame_flag),
	.D(n85),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Address_seq_reg[0]  (
	.SI(test_si),
	.SE(n111),
	.RN(FE_OFN3_O_RST2),
	.Q(Address_seq[0]),
	.D(n84),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Address_seq_reg[1]  (
	.SI(Address_seq[0]),
	.SE(n112),
	.RN(FE_OFN3_O_RST2),
	.Q(Address_seq[1]),
	.D(n83),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Address_seq_reg[3]  (
	.SI(Address_seq[2]),
	.SE(n108),
	.RN(FE_OFN3_O_RST2),
	.Q(Address_seq[3]),
	.D(n81),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Address_seq_reg[2]  (
	.SI(Address_seq[1]),
	.SE(n113),
	.RN(FE_OFN3_O_RST2),
	.Q(Address_seq[2]),
	.D(n82),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U133 (
	.Y(n105),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U135 (
	.Y(n107),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U136 (
	.Y(n108),
	.A(n111), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U137 (
	.Y(n109),
	.A(n112), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U138 (
	.Y(n110),
	.A(n113), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U139 (
	.Y(n111),
	.A(n107), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U140 (
	.Y(n112),
	.A(n107), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U141 (
	.Y(n113),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U142 (
	.Y(n114),
	.A(ALU_OUT_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(clk_div_en),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Reg_File_ADD_WIDTH4_RdWr_WIDTH8_RegF_DEPTH16_test_1 (
	RdEn, 
	WrEn, 
	CLK, 
	RST, 
	ADDRESS, 
	Wr_DATA, 
	Rd_DATA, 
	Rd_DATA_VLD, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si2, 
	test_si1, 
	test_so1, 
	test_se, 
	FE_OFN0_O_RST2, 
	FE_OFN2_O_RST2, 
	FE_OFN3_O_RST2, 
	O_CLK1__L5_N1, 
	O_CLK1__L5_N2, 
	O_CLK1__L5_N3, 
	O_CLK1__L5_N4, 
	O_CLK1__L5_N5, 
	O_CLK1__L5_N7, 
	VDD, 
	VSS);
   input RdEn;
   input WrEn;
   input CLK;
   input RST;
   input [3:0] ADDRESS;
   input [7:0] Wr_DATA;
   output [7:0] Rd_DATA;
   output Rd_DATA_VLD;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si2;
   input test_si1;
   output test_so1;
   input test_se;
   input FE_OFN0_O_RST2;
   input FE_OFN2_O_RST2;
   input FE_OFN3_O_RST2;
   input O_CLK1__L5_N1;
   input O_CLK1__L5_N2;
   input O_CLK1__L5_N3;
   input O_CLK1__L5_N4;
   input O_CLK1__L5_N5;
   input O_CLK1__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire FE_OFN1_O_RST2;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire n275;
   wire n466;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire \REG_FILE[4][7] ;
   wire \REG_FILE[4][6] ;
   wire \REG_FILE[4][5] ;
   wire \REG_FILE[4][4] ;
   wire \REG_FILE[4][3] ;
   wire \REG_FILE[4][2] ;
   wire \REG_FILE[4][1] ;
   wire \REG_FILE[4][0] ;
   wire \REG_FILE[5][7] ;
   wire \REG_FILE[5][6] ;
   wire \REG_FILE[5][5] ;
   wire \REG_FILE[5][4] ;
   wire \REG_FILE[5][3] ;
   wire \REG_FILE[5][2] ;
   wire \REG_FILE[5][1] ;
   wire \REG_FILE[5][0] ;
   wire \REG_FILE[6][7] ;
   wire \REG_FILE[6][6] ;
   wire \REG_FILE[6][5] ;
   wire \REG_FILE[6][4] ;
   wire \REG_FILE[6][3] ;
   wire \REG_FILE[6][2] ;
   wire \REG_FILE[6][1] ;
   wire \REG_FILE[6][0] ;
   wire \REG_FILE[7][7] ;
   wire \REG_FILE[7][6] ;
   wire \REG_FILE[7][5] ;
   wire \REG_FILE[7][4] ;
   wire \REG_FILE[7][3] ;
   wire \REG_FILE[7][2] ;
   wire \REG_FILE[7][1] ;
   wire \REG_FILE[7][0] ;
   wire \REG_FILE[8][7] ;
   wire \REG_FILE[8][6] ;
   wire \REG_FILE[8][5] ;
   wire \REG_FILE[8][4] ;
   wire \REG_FILE[8][3] ;
   wire \REG_FILE[8][2] ;
   wire \REG_FILE[8][1] ;
   wire \REG_FILE[8][0] ;
   wire \REG_FILE[9][7] ;
   wire \REG_FILE[9][6] ;
   wire \REG_FILE[9][5] ;
   wire \REG_FILE[9][4] ;
   wire \REG_FILE[9][3] ;
   wire \REG_FILE[9][2] ;
   wire \REG_FILE[9][1] ;
   wire \REG_FILE[9][0] ;
   wire \REG_FILE[10][7] ;
   wire \REG_FILE[10][6] ;
   wire \REG_FILE[10][5] ;
   wire \REG_FILE[10][4] ;
   wire \REG_FILE[10][3] ;
   wire \REG_FILE[10][2] ;
   wire \REG_FILE[10][1] ;
   wire \REG_FILE[10][0] ;
   wire \REG_FILE[11][7] ;
   wire \REG_FILE[11][6] ;
   wire \REG_FILE[11][5] ;
   wire \REG_FILE[11][4] ;
   wire \REG_FILE[11][3] ;
   wire \REG_FILE[11][2] ;
   wire \REG_FILE[11][1] ;
   wire \REG_FILE[11][0] ;
   wire \REG_FILE[12][7] ;
   wire \REG_FILE[12][6] ;
   wire \REG_FILE[12][5] ;
   wire \REG_FILE[12][4] ;
   wire \REG_FILE[12][3] ;
   wire \REG_FILE[12][2] ;
   wire \REG_FILE[12][1] ;
   wire \REG_FILE[12][0] ;
   wire \REG_FILE[13][7] ;
   wire \REG_FILE[13][6] ;
   wire \REG_FILE[13][5] ;
   wire \REG_FILE[13][4] ;
   wire \REG_FILE[13][3] ;
   wire \REG_FILE[13][2] ;
   wire \REG_FILE[13][1] ;
   wire \REG_FILE[13][0] ;
   wire \REG_FILE[14][7] ;
   wire \REG_FILE[14][6] ;
   wire \REG_FILE[14][5] ;
   wire \REG_FILE[14][4] ;
   wire \REG_FILE[14][3] ;
   wire \REG_FILE[14][2] ;
   wire \REG_FILE[14][1] ;
   wire \REG_FILE[14][0] ;
   wire \REG_FILE[15][7] ;
   wire \REG_FILE[15][6] ;
   wire \REG_FILE[15][5] ;
   wire \REG_FILE[15][4] ;
   wire \REG_FILE[15][3] ;
   wire \REG_FILE[15][2] ;
   wire \REG_FILE[15][1] ;
   wire \REG_FILE[15][0] ;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n1;
   wire n3;
   wire n12;
   wire n13;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n436;
   wire n2;

   assign N11 = ADDRESS[0] ;
   assign N12 = ADDRESS[1] ;
   assign N13 = ADDRESS[2] ;
   assign N14 = ADDRESS[3] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M FE_OFC1_O_RST2 (
	.Y(FE_OFN1_O_RST2),
	.A(FE_OFN0_O_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U3 (
	.Y(n1),
	.A(n275), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U4 (
	.Y(REG1[1]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U7 (
	.Y(REG2[7]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U15 (
	.Y(n264),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(n22),
	.B(n249),
	.A(n264), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(n17),
	.B(n250),
	.A(n264), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(n32),
	.B(n247),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U19 (
	.Y(n34),
	.B(n248),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U20 (
	.Y(n20),
	.B(n248),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U21 (
	.Y(n18),
	.B(n247),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n250),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(n28),
	.B(N13),
	.A(n249), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U25 (
	.Y(n25),
	.B(N13),
	.A(n250), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U26 (
	.Y(n180),
	.S1(n249),
	.S0(n247),
	.D(REG3[0]),
	.C(REG2[0]),
	.B(REG1[0]),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U27 (
	.Y(n188),
	.S1(n249),
	.S0(n247),
	.D(n476),
	.C(REG2[2]),
	.B(REG1[2]),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U28 (
	.Y(n196),
	.S1(n249),
	.S0(n247),
	.D(n474),
	.C(REG2[4]),
	.B(REG1[4]),
	.A(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U29 (
	.Y(n200),
	.S1(n249),
	.S0(n247),
	.D(REG3[5]),
	.C(REG2[5]),
	.B(REG1[5]),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U30 (
	.Y(n204),
	.S1(n249),
	.S0(n247),
	.D(n473),
	.C(REG2[6]),
	.B(REG1[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U31 (
	.Y(n208),
	.S1(n249),
	.S0(n247),
	.D(n472),
	.C(REG2[7]),
	.B(REG1[7]),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U32 (
	.Y(n184),
	.S1(n249),
	.S0(n247),
	.D(n477),
	.C(REG2[1]),
	.B(REG1[1]),
	.A(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U33 (
	.Y(n267),
	.A(Wr_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U64 (
	.Y(n16),
	.B(n18),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U65 (
	.Y(n21),
	.B(n18),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U66 (
	.Y(n23),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U75 (
	.Y(n19),
	.B(n17),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U76 (
	.Y(n31),
	.B(n17),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U77 (
	.Y(n33),
	.B(n17),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U78 (
	.Y(n35),
	.B(n22),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U79 (
	.Y(n36),
	.B(n22),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U88 (
	.Y(n265),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U91 (
	.Y(n37),
	.B(n25),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U92 (
	.Y(n38),
	.B(n25),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U93 (
	.Y(n39),
	.B(n28),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U94 (
	.Y(n41),
	.B(n28),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U95 (
	.Y(n24),
	.B(n18),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U96 (
	.Y(n26),
	.B(n20),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U97 (
	.Y(n27),
	.B(n18),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U98 (
	.Y(n30),
	.B(n20),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U99 (
	.Y(n249),
	.A(n250), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX6M U100 (
	.Y(n247),
	.A(n248), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U101 (
	.Y(n14),
	.B(RdEn),
	.A(n266), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U102 (
	.Y(n266),
	.A(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U103 (
	.Y(n15),
	.B(n266),
	.A(RdEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U104 (
	.Y(n40),
	.B(N14),
	.AN(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U105 (
	.Y(n29),
	.B(n14),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n248),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U107 (
	.Y(n274),
	.A(Wr_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U108 (
	.Y(n273),
	.A(Wr_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U109 (
	.Y(n272),
	.A(Wr_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U110 (
	.Y(n271),
	.A(Wr_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U111 (
	.Y(n270),
	.A(Wr_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U112 (
	.Y(n269),
	.A(Wr_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U113 (
	.Y(n268),
	.A(Wr_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U115 (
	.Y(n51),
	.B1(n274),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U116 (
	.Y(n52),
	.B1(n273),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U117 (
	.Y(n53),
	.B1(n272),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n54),
	.B1(n271),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n55),
	.B1(n270),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n56),
	.B1(n269),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n57),
	.B1(n268),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n59),
	.B1(n19),
	.B0(n274),
	.A1N(n19),
	.A0N(\REG_FILE[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n60),
	.B1(n19),
	.B0(n273),
	.A1N(n19),
	.A0N(\REG_FILE[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n61),
	.B1(n19),
	.B0(n272),
	.A1N(n19),
	.A0N(\REG_FILE[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U125 (
	.Y(n62),
	.B1(n19),
	.B0(n271),
	.A1N(n19),
	.A0N(\REG_FILE[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U126 (
	.Y(n63),
	.B1(n19),
	.B0(n270),
	.A1N(n19),
	.A0N(\REG_FILE[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U127 (
	.Y(n64),
	.B1(n19),
	.B0(n269),
	.A1N(n19),
	.A0N(\REG_FILE[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U128 (
	.Y(n65),
	.B1(n19),
	.B0(n268),
	.A1N(n19),
	.A0N(\REG_FILE[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U129 (
	.Y(n67),
	.B1(n21),
	.B0(n274),
	.A1N(n21),
	.A0N(\REG_FILE[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U130 (
	.Y(n68),
	.B1(n21),
	.B0(n273),
	.A1N(n21),
	.A0N(\REG_FILE[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U131 (
	.Y(n69),
	.B1(n21),
	.B0(n272),
	.A1N(n21),
	.A0N(\REG_FILE[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U132 (
	.Y(n70),
	.B1(n21),
	.B0(n271),
	.A1N(n21),
	.A0N(\REG_FILE[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U133 (
	.Y(n71),
	.B1(n21),
	.B0(n270),
	.A1N(n21),
	.A0N(\REG_FILE[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U134 (
	.Y(n72),
	.B1(n21),
	.B0(n269),
	.A1N(n21),
	.A0N(\REG_FILE[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U135 (
	.Y(n73),
	.B1(n21),
	.B0(n268),
	.A1N(n21),
	.A0N(\REG_FILE[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n75),
	.B1(n23),
	.B0(n274),
	.A1N(n23),
	.A0N(\REG_FILE[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n76),
	.B1(n23),
	.B0(n273),
	.A1N(n23),
	.A0N(\REG_FILE[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n77),
	.B1(n23),
	.B0(n272),
	.A1N(n23),
	.A0N(\REG_FILE[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n78),
	.B1(n23),
	.B0(n271),
	.A1N(n23),
	.A0N(\REG_FILE[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n79),
	.B1(n23),
	.B0(n270),
	.A1N(n23),
	.A0N(\REG_FILE[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n80),
	.B1(n23),
	.B0(n269),
	.A1N(n23),
	.A0N(\REG_FILE[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n81),
	.B1(n23),
	.B0(n268),
	.A1N(n23),
	.A0N(\REG_FILE[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n83),
	.B1(n24),
	.B0(n274),
	.A1N(n24),
	.A0N(\REG_FILE[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n84),
	.B1(n24),
	.B0(n273),
	.A1N(n24),
	.A0N(\REG_FILE[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n85),
	.B1(n24),
	.B0(n272),
	.A1N(n24),
	.A0N(\REG_FILE[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n86),
	.B1(n24),
	.B0(n271),
	.A1N(n24),
	.A0N(\REG_FILE[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n87),
	.B1(n24),
	.B0(n270),
	.A1N(n24),
	.A0N(\REG_FILE[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n88),
	.B1(n24),
	.B0(n269),
	.A1N(n24),
	.A0N(\REG_FILE[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U149 (
	.Y(n89),
	.B1(n24),
	.B0(n268),
	.A1N(n24),
	.A0N(\REG_FILE[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U150 (
	.Y(n91),
	.B1(n26),
	.B0(n274),
	.A1N(n26),
	.A0N(\REG_FILE[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U151 (
	.Y(n92),
	.B1(n26),
	.B0(n273),
	.A1N(n26),
	.A0N(\REG_FILE[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U152 (
	.Y(n93),
	.B1(n26),
	.B0(n272),
	.A1N(n26),
	.A0N(\REG_FILE[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U153 (
	.Y(n94),
	.B1(n26),
	.B0(n271),
	.A1N(n26),
	.A0N(\REG_FILE[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U154 (
	.Y(n95),
	.B1(n26),
	.B0(n270),
	.A1N(n26),
	.A0N(\REG_FILE[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U155 (
	.Y(n96),
	.B1(n26),
	.B0(n269),
	.A1N(n26),
	.A0N(\REG_FILE[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U156 (
	.Y(n97),
	.B1(n26),
	.B0(n268),
	.A1N(n26),
	.A0N(\REG_FILE[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U157 (
	.Y(n99),
	.B1(n27),
	.B0(n274),
	.A1N(n27),
	.A0N(\REG_FILE[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U158 (
	.Y(n100),
	.B1(n27),
	.B0(n273),
	.A1N(n27),
	.A0N(\REG_FILE[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U159 (
	.Y(n101),
	.B1(n27),
	.B0(n272),
	.A1N(n27),
	.A0N(\REG_FILE[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U160 (
	.Y(n102),
	.B1(n27),
	.B0(n271),
	.A1N(n27),
	.A0N(\REG_FILE[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U161 (
	.Y(n103),
	.B1(n27),
	.B0(n270),
	.A1N(n27),
	.A0N(\REG_FILE[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U162 (
	.Y(n104),
	.B1(n27),
	.B0(n269),
	.A1N(n27),
	.A0N(\REG_FILE[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U163 (
	.Y(n105),
	.B1(n27),
	.B0(n268),
	.A1N(n27),
	.A0N(\REG_FILE[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U164 (
	.Y(n107),
	.B1(n30),
	.B0(n274),
	.A1N(n30),
	.A0N(\REG_FILE[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U165 (
	.Y(n108),
	.B1(n30),
	.B0(n273),
	.A1N(n30),
	.A0N(\REG_FILE[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U166 (
	.Y(n109),
	.B1(n30),
	.B0(n272),
	.A1N(n30),
	.A0N(\REG_FILE[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U167 (
	.Y(n110),
	.B1(n30),
	.B0(n271),
	.A1N(n30),
	.A0N(test_so1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U168 (
	.Y(n111),
	.B1(n30),
	.B0(n270),
	.A1N(n30),
	.A0N(\REG_FILE[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U169 (
	.Y(n112),
	.B1(n30),
	.B0(n269),
	.A1N(n30),
	.A0N(\REG_FILE[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U170 (
	.Y(n113),
	.B1(n30),
	.B0(n268),
	.A1N(n30),
	.A0N(\REG_FILE[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U171 (
	.Y(n115),
	.B1(n31),
	.B0(n274),
	.A1N(n31),
	.A0N(\REG_FILE[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U172 (
	.Y(n116),
	.B1(n31),
	.B0(n273),
	.A1N(n31),
	.A0N(\REG_FILE[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U173 (
	.Y(n117),
	.B1(n31),
	.B0(n272),
	.A1N(n31),
	.A0N(\REG_FILE[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U174 (
	.Y(n118),
	.B1(n31),
	.B0(n271),
	.A1N(n31),
	.A0N(\REG_FILE[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U175 (
	.Y(n119),
	.B1(n31),
	.B0(n270),
	.A1N(n31),
	.A0N(\REG_FILE[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U176 (
	.Y(n120),
	.B1(n31),
	.B0(n269),
	.A1N(n31),
	.A0N(\REG_FILE[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U177 (
	.Y(n121),
	.B1(n31),
	.B0(n268),
	.A1N(n31),
	.A0N(\REG_FILE[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U178 (
	.Y(n123),
	.B1(n33),
	.B0(n274),
	.A1N(n33),
	.A0N(\REG_FILE[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U179 (
	.Y(n124),
	.B1(n33),
	.B0(n273),
	.A1N(n33),
	.A0N(\REG_FILE[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U180 (
	.Y(n125),
	.B1(n33),
	.B0(n272),
	.A1N(n33),
	.A0N(\REG_FILE[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U181 (
	.Y(n126),
	.B1(n33),
	.B0(n271),
	.A1N(n33),
	.A0N(\REG_FILE[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U182 (
	.Y(n127),
	.B1(n33),
	.B0(n270),
	.A1N(n33),
	.A0N(\REG_FILE[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U183 (
	.Y(n128),
	.B1(n33),
	.B0(n269),
	.A1N(n33),
	.A0N(\REG_FILE[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U184 (
	.Y(n129),
	.B1(n33),
	.B0(n268),
	.A1N(n33),
	.A0N(\REG_FILE[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U185 (
	.Y(n131),
	.B1(n35),
	.B0(n274),
	.A1N(n35),
	.A0N(\REG_FILE[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U186 (
	.Y(n132),
	.B1(n35),
	.B0(n273),
	.A1N(n35),
	.A0N(\REG_FILE[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U187 (
	.Y(n133),
	.B1(n35),
	.B0(n272),
	.A1N(n35),
	.A0N(\REG_FILE[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U188 (
	.Y(n134),
	.B1(n35),
	.B0(n271),
	.A1N(n35),
	.A0N(\REG_FILE[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U189 (
	.Y(n135),
	.B1(n35),
	.B0(n270),
	.A1N(n35),
	.A0N(\REG_FILE[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U190 (
	.Y(n136),
	.B1(n35),
	.B0(n269),
	.A1N(n35),
	.A0N(\REG_FILE[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U191 (
	.Y(n137),
	.B1(n35),
	.B0(n268),
	.A1N(n35),
	.A0N(\REG_FILE[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U192 (
	.Y(n139),
	.B1(n36),
	.B0(n274),
	.A1N(n36),
	.A0N(\REG_FILE[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U193 (
	.Y(n140),
	.B1(n36),
	.B0(n273),
	.A1N(n36),
	.A0N(\REG_FILE[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U194 (
	.Y(n141),
	.B1(n36),
	.B0(n272),
	.A1N(n36),
	.A0N(\REG_FILE[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U195 (
	.Y(n142),
	.B1(n36),
	.B0(n271),
	.A1N(n36),
	.A0N(\REG_FILE[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U196 (
	.Y(n143),
	.B1(n36),
	.B0(n270),
	.A1N(n36),
	.A0N(\REG_FILE[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U197 (
	.Y(n144),
	.B1(n36),
	.B0(n269),
	.A1N(n36),
	.A0N(\REG_FILE[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U198 (
	.Y(n145),
	.B1(n36),
	.B0(n268),
	.A1N(n36),
	.A0N(\REG_FILE[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U199 (
	.Y(n147),
	.B1(n37),
	.B0(n274),
	.A1N(n37),
	.A0N(REG3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U200 (
	.Y(n148),
	.B1(n37),
	.B0(n273),
	.A1N(n37),
	.A0N(n477), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U201 (
	.Y(n149),
	.B1(n37),
	.B0(n272),
	.A1N(n37),
	.A0N(n476), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U202 (
	.Y(n150),
	.B1(n37),
	.B0(n271),
	.A1N(n37),
	.A0N(n475), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U203 (
	.Y(n151),
	.B1(n37),
	.B0(n270),
	.A1N(n37),
	.A0N(n474), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U204 (
	.Y(n153),
	.B1(n37),
	.B0(n268),
	.A1N(n37),
	.A0N(n473), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U205 (
	.Y(n156),
	.B1(n38),
	.B0(n273),
	.A1N(n38),
	.A0N(REG2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U206 (
	.Y(n157),
	.B1(n38),
	.B0(n272),
	.A1N(n38),
	.A0N(REG2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n158),
	.B1(n38),
	.B0(n271),
	.A1N(n38),
	.A0N(REG2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n159),
	.B1(n38),
	.B0(n270),
	.A1N(n38),
	.A0N(REG2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n160),
	.B1(n38),
	.B0(n269),
	.A1N(n38),
	.A0N(REG2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n161),
	.B1(n38),
	.B0(n268),
	.A1N(n38),
	.A0N(REG2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n163),
	.B1(n39),
	.B0(n274),
	.A1N(n39),
	.A0N(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n164),
	.B1(n39),
	.B0(n273),
	.A1N(n39),
	.A0N(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n165),
	.B1(n39),
	.B0(n272),
	.A1N(n39),
	.A0N(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n166),
	.B1(n39),
	.B0(n271),
	.A1N(n39),
	.A0N(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n167),
	.B1(n39),
	.B0(n270),
	.A1N(n39),
	.A0N(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n168),
	.B1(n39),
	.B0(n269),
	.A1N(n39),
	.A0N(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n169),
	.B1(n39),
	.B0(n268),
	.A1N(n39),
	.A0N(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n171),
	.B1(n41),
	.B0(n274),
	.A1N(n41),
	.A0N(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n172),
	.B1(n41),
	.B0(n273),
	.A1N(n41),
	.A0N(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n173),
	.B1(n41),
	.B0(n272),
	.A1N(n41),
	.A0N(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n174),
	.B1(n41),
	.B0(n271),
	.A1N(n41),
	.A0N(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n175),
	.B1(n41),
	.B0(n270),
	.A1N(n41),
	.A0N(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n176),
	.B1(n41),
	.B0(n269),
	.A1N(n41),
	.A0N(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n177),
	.B1(n41),
	.B0(n268),
	.A1N(n41),
	.A0N(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n58),
	.B1(n267),
	.B0(n16),
	.A1N(n16),
	.A0N(\REG_FILE[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n66),
	.B1(n19),
	.B0(n267),
	.A1N(n19),
	.A0N(\REG_FILE[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n74),
	.B1(n21),
	.B0(n267),
	.A1N(n21),
	.A0N(\REG_FILE[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n82),
	.B1(n23),
	.B0(n267),
	.A1N(n23),
	.A0N(\REG_FILE[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n90),
	.B1(n24),
	.B0(n267),
	.A1N(n24),
	.A0N(\REG_FILE[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n98),
	.B1(n26),
	.B0(n267),
	.A1N(n26),
	.A0N(\REG_FILE[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n106),
	.B1(n27),
	.B0(n267),
	.A1N(n27),
	.A0N(\REG_FILE[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n114),
	.B1(n30),
	.B0(n267),
	.A1N(n30),
	.A0N(\REG_FILE[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n122),
	.B1(n31),
	.B0(n267),
	.A1N(n31),
	.A0N(\REG_FILE[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n130),
	.B1(n33),
	.B0(n267),
	.A1N(n33),
	.A0N(\REG_FILE[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n138),
	.B1(n35),
	.B0(n267),
	.A1N(n35),
	.A0N(\REG_FILE[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n146),
	.B1(n36),
	.B0(n267),
	.A1N(n36),
	.A0N(\REG_FILE[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n154),
	.B1(n37),
	.B0(n267),
	.A1N(n37),
	.A0N(n472), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U238 (
	.Y(n170),
	.B1(n39),
	.B0(n267),
	.A1N(n39),
	.A0N(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n178),
	.B1(n41),
	.B0(n267),
	.A1N(n41),
	.A0N(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U240 (
	.Y(n152),
	.B1(n37),
	.B0(n269),
	.A1N(n37),
	.A0N(REG3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U241 (
	.Y(n155),
	.B1(n38),
	.B0(n274),
	.A1N(n38),
	.A0N(REG2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U242 (
	.Y(n162),
	.B1(n38),
	.B0(n267),
	.A1N(n38),
	.A0N(REG2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U243 (
	.Y(n187),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][2] ),
	.C(\REG_FILE[6][2] ),
	.B(\REG_FILE[5][2] ),
	.A(\REG_FILE[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U244 (
	.Y(n191),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][3] ),
	.C(\REG_FILE[6][3] ),
	.B(\REG_FILE[5][3] ),
	.A(\REG_FILE[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U245 (
	.Y(n195),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][4] ),
	.C(\REG_FILE[6][4] ),
	.B(\REG_FILE[5][4] ),
	.A(\REG_FILE[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U246 (
	.Y(n199),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][5] ),
	.C(\REG_FILE[6][5] ),
	.B(\REG_FILE[5][5] ),
	.A(\REG_FILE[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U247 (
	.Y(n203),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][6] ),
	.C(\REG_FILE[6][6] ),
	.B(\REG_FILE[5][6] ),
	.A(\REG_FILE[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U248 (
	.Y(n207),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][7] ),
	.C(\REG_FILE[6][7] ),
	.B(\REG_FILE[5][7] ),
	.A(\REG_FILE[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U249 (
	.Y(n185),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][2] ),
	.C(\REG_FILE[14][2] ),
	.B(\REG_FILE[13][2] ),
	.A(\REG_FILE[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U250 (
	.Y(n189),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][3] ),
	.C(\REG_FILE[14][3] ),
	.B(\REG_FILE[13][3] ),
	.A(\REG_FILE[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U251 (
	.Y(n193),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][4] ),
	.C(\REG_FILE[14][4] ),
	.B(\REG_FILE[13][4] ),
	.A(\REG_FILE[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U252 (
	.Y(n197),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][5] ),
	.C(\REG_FILE[14][5] ),
	.B(\REG_FILE[13][5] ),
	.A(\REG_FILE[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U253 (
	.Y(n201),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][6] ),
	.C(\REG_FILE[14][6] ),
	.B(\REG_FILE[13][6] ),
	.A(\REG_FILE[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U254 (
	.Y(n205),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][7] ),
	.C(\REG_FILE[14][7] ),
	.B(\REG_FILE[13][7] ),
	.A(\REG_FILE[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U255 (
	.Y(n183),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[7][1] ),
	.C(\REG_FILE[6][1] ),
	.B(\REG_FILE[5][1] ),
	.A(\REG_FILE[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U256 (
	.Y(n44),
	.B1(n15),
	.B0(Rd_DATA[1]),
	.A1(n265),
	.A0(N42), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U257 (
	.Y(N42),
	.S1(N13),
	.S0(N14),
	.D(n181),
	.C(n183),
	.B(n182),
	.A(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U258 (
	.Y(n182),
	.S1(N12),
	.S0(N11),
	.D(\REG_FILE[11][1] ),
	.C(\REG_FILE[10][1] ),
	.B(\REG_FILE[9][1] ),
	.A(\REG_FILE[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U259 (
	.Y(n181),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][1] ),
	.C(\REG_FILE[14][1] ),
	.B(\REG_FILE[13][1] ),
	.A(\REG_FILE[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U260 (
	.Y(n45),
	.B1(n15),
	.B0(Rd_DATA[2]),
	.A1(n265),
	.A0(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U261 (
	.Y(N41),
	.S1(N13),
	.S0(N14),
	.D(n185),
	.C(n187),
	.B(n186),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U262 (
	.Y(n186),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[11][2] ),
	.C(\REG_FILE[10][2] ),
	.B(\REG_FILE[9][2] ),
	.A(\REG_FILE[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U263 (
	.Y(n46),
	.B1(n15),
	.B0(Rd_DATA[3]),
	.A1(n265),
	.A0(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U264 (
	.Y(N40),
	.S1(N13),
	.S0(N14),
	.D(n189),
	.C(n191),
	.B(n190),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U265 (
	.Y(n192),
	.S1(n249),
	.S0(n247),
	.D(n475),
	.C(REG2[3]),
	.B(REG1[3]),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U266 (
	.Y(n190),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[11][3] ),
	.C(\REG_FILE[10][3] ),
	.B(\REG_FILE[9][3] ),
	.A(test_so1), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U267 (
	.Y(n47),
	.B1(n15),
	.B0(Rd_DATA[4]),
	.A1(n265),
	.A0(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U268 (
	.Y(N39),
	.S1(N13),
	.S0(N14),
	.D(n193),
	.C(n195),
	.B(n194),
	.A(n196), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U269 (
	.Y(n194),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[11][4] ),
	.C(\REG_FILE[10][4] ),
	.B(\REG_FILE[9][4] ),
	.A(\REG_FILE[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U270 (
	.Y(n48),
	.B1(n15),
	.B0(Rd_DATA[5]),
	.A1(n265),
	.A0(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U271 (
	.Y(N38),
	.S1(N13),
	.S0(N14),
	.D(n197),
	.C(n199),
	.B(n198),
	.A(n200), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U272 (
	.Y(n198),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[11][5] ),
	.C(\REG_FILE[10][5] ),
	.B(\REG_FILE[9][5] ),
	.A(\REG_FILE[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U273 (
	.Y(n49),
	.B1(n15),
	.B0(Rd_DATA[6]),
	.A1(n265),
	.A0(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U274 (
	.Y(N37),
	.S1(N13),
	.S0(N14),
	.D(n201),
	.C(n203),
	.B(n202),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U275 (
	.Y(n202),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[11][6] ),
	.C(\REG_FILE[10][6] ),
	.B(\REG_FILE[9][6] ),
	.A(\REG_FILE[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U276 (
	.Y(n50),
	.B1(n15),
	.B0(Rd_DATA[7]),
	.A1(n265),
	.A0(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U277 (
	.Y(N36),
	.S1(N13),
	.S0(N14),
	.D(n205),
	.C(n207),
	.B(n206),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U278 (
	.Y(n206),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[11][7] ),
	.C(\REG_FILE[10][7] ),
	.B(\REG_FILE[9][7] ),
	.A(\REG_FILE[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U279 (
	.Y(n179),
	.S1(n249),
	.S0(N11),
	.D(\REG_FILE[7][0] ),
	.C(\REG_FILE[6][0] ),
	.B(\REG_FILE[5][0] ),
	.A(\REG_FILE[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U280 (
	.Y(n12),
	.S1(n249),
	.S0(n247),
	.D(\REG_FILE[15][0] ),
	.C(\REG_FILE[14][0] ),
	.B(\REG_FILE[13][0] ),
	.A(\REG_FILE[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U281 (
	.Y(n43),
	.B1(n15),
	.B0(Rd_DATA[0]),
	.A1(n265),
	.A0(N43), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U282 (
	.Y(N43),
	.S1(N13),
	.S0(N14),
	.D(n12),
	.C(n179),
	.B(n13),
	.A(n180), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U283 (
	.Y(n13),
	.S1(N12),
	.S0(N11),
	.D(\REG_FILE[11][0] ),
	.C(\REG_FILE[10][0] ),
	.B(\REG_FILE[9][0] ),
	.A(\REG_FILE[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U284 (
	.Y(n42),
	.B0(n265),
	.A1(n14),
	.A0(Rd_DATA_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \REG_FILE_reg[1][0]  (
	.SI(REG0[7]),
	.SE(n301),
	.RN(FE_OFN3_O_RST2),
	.Q(n466),
	.D(n163),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \REG_FILE_reg[2][5]  (
	.SI(REG2[4]),
	.SE(n296),
	.RN(FE_OFN3_O_RST2),
	.Q(REG2[5]),
	.D(n160),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][7]  (
	.SI(\REG_FILE[5][6] ),
	.SE(n424),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][7] ),
	.D(n138),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][6]  (
	.SI(\REG_FILE[5][5] ),
	.SE(n361),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][6] ),
	.D(n137),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][5]  (
	.SI(\REG_FILE[5][4] ),
	.SE(n423),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][5] ),
	.D(n136),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][4]  (
	.SI(\REG_FILE[5][3] ),
	.SE(n360),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][4] ),
	.D(n135),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][3]  (
	.SI(\REG_FILE[5][2] ),
	.SE(n422),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][3] ),
	.D(n134),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][2]  (
	.SI(\REG_FILE[5][1] ),
	.SE(n359),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][2] ),
	.D(n133),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][1]  (
	.SI(\REG_FILE[5][0] ),
	.SE(n421),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][1] ),
	.D(n132),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[5][0]  (
	.SI(\REG_FILE[4][7] ),
	.SE(n358),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[5][0] ),
	.D(n131),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][7]  (
	.SI(\REG_FILE[9][6] ),
	.SE(n285),
	.RN(RST),
	.Q(\REG_FILE[9][7] ),
	.D(n106),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][6]  (
	.SI(\REG_FILE[9][5] ),
	.SE(n286),
	.RN(RST),
	.Q(\REG_FILE[9][6] ),
	.D(n105),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][5]  (
	.SI(\REG_FILE[9][4] ),
	.SE(n305),
	.RN(RST),
	.Q(\REG_FILE[9][5] ),
	.D(n104),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][4]  (
	.SI(\REG_FILE[9][3] ),
	.SE(n377),
	.RN(RST),
	.Q(\REG_FILE[9][4] ),
	.D(n103),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][3]  (
	.SI(\REG_FILE[9][2] ),
	.SE(n376),
	.RN(RST),
	.Q(\REG_FILE[9][3] ),
	.D(n102),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][2]  (
	.SI(\REG_FILE[9][1] ),
	.SE(n314),
	.RN(RST),
	.Q(\REG_FILE[9][2] ),
	.D(n101),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][1]  (
	.SI(\REG_FILE[9][0] ),
	.SE(n287),
	.RN(RST),
	.Q(\REG_FILE[9][1] ),
	.D(n100),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[9][0]  (
	.SI(\REG_FILE[8][7] ),
	.SE(n288),
	.RN(RST),
	.Q(\REG_FILE[9][0] ),
	.D(n99),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][7]  (
	.SI(\REG_FILE[13][6] ),
	.SE(n330),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][7] ),
	.D(n74),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][6]  (
	.SI(\REG_FILE[13][5] ),
	.SE(n392),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][6] ),
	.D(n73),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][5]  (
	.SI(\REG_FILE[13][4] ),
	.SE(n329),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][5] ),
	.D(n72),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][4]  (
	.SI(\REG_FILE[13][3] ),
	.SE(n391),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][4] ),
	.D(n71),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][3]  (
	.SI(\REG_FILE[13][2] ),
	.SE(n328),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][3] ),
	.D(n70),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][2]  (
	.SI(\REG_FILE[13][1] ),
	.SE(n390),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][2] ),
	.D(n69),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][1]  (
	.SI(\REG_FILE[13][0] ),
	.SE(n327),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][1] ),
	.D(n68),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[13][0]  (
	.SI(\REG_FILE[12][7] ),
	.SE(n389),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[13][0] ),
	.D(n67),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][7]  (
	.SI(\REG_FILE[7][6] ),
	.SE(n432),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][7] ),
	.D(n122),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][6]  (
	.SI(\REG_FILE[7][5] ),
	.SE(n369),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][6] ),
	.D(n121),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][5]  (
	.SI(\REG_FILE[7][4] ),
	.SE(n431),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][5] ),
	.D(n120),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][4]  (
	.SI(\REG_FILE[7][3] ),
	.SE(n368),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][4] ),
	.D(n119),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][3]  (
	.SI(\REG_FILE[7][2] ),
	.SE(n430),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][3] ),
	.D(n118),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][2]  (
	.SI(\REG_FILE[7][1] ),
	.SE(n367),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][2] ),
	.D(n117),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][1]  (
	.SI(\REG_FILE[7][0] ),
	.SE(n429),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][1] ),
	.D(n116),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[7][0]  (
	.SI(\REG_FILE[6][7] ),
	.SE(n366),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[7][0] ),
	.D(n115),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][7]  (
	.SI(\REG_FILE[11][6] ),
	.SE(n322),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][7] ),
	.D(n90),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][6]  (
	.SI(\REG_FILE[11][5] ),
	.SE(n384),
	.RN(RST),
	.Q(\REG_FILE[11][6] ),
	.D(n89),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][5]  (
	.SI(\REG_FILE[11][4] ),
	.SE(n321),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][5] ),
	.D(n88),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][4]  (
	.SI(\REG_FILE[11][3] ),
	.SE(n383),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][4] ),
	.D(n87),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][3]  (
	.SI(\REG_FILE[11][2] ),
	.SE(n320),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][3] ),
	.D(n86),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][2]  (
	.SI(\REG_FILE[11][1] ),
	.SE(n382),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][2] ),
	.D(n85),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][1]  (
	.SI(\REG_FILE[11][0] ),
	.SE(n319),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][1] ),
	.D(n84),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[11][0]  (
	.SI(\REG_FILE[10][7] ),
	.SE(n381),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[11][0] ),
	.D(n83),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][7]  (
	.SI(\REG_FILE[15][6] ),
	.SE(n338),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[15][7] ),
	.D(n58),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][6]  (
	.SI(\REG_FILE[15][5] ),
	.SE(n400),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[15][6] ),
	.D(n57),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][5]  (
	.SI(\REG_FILE[15][4] ),
	.SE(n337),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[15][5] ),
	.D(n56),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][4]  (
	.SI(\REG_FILE[15][3] ),
	.SE(n399),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[15][4] ),
	.D(n55),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][3]  (
	.SI(\REG_FILE[15][2] ),
	.SE(n336),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[15][3] ),
	.D(n54),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][2]  (
	.SI(\REG_FILE[15][1] ),
	.SE(n398),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[15][2] ),
	.D(n53),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][1]  (
	.SI(\REG_FILE[15][0] ),
	.SE(n335),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[15][1] ),
	.D(n52),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[15][0]  (
	.SI(\REG_FILE[14][7] ),
	.SE(n397),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[15][0] ),
	.D(n51),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][7]  (
	.SI(\REG_FILE[6][6] ),
	.SE(n428),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][7] ),
	.D(n130),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][6]  (
	.SI(\REG_FILE[6][5] ),
	.SE(n365),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][6] ),
	.D(n129),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][5]  (
	.SI(\REG_FILE[6][4] ),
	.SE(n427),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][5] ),
	.D(n128),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][4]  (
	.SI(\REG_FILE[6][3] ),
	.SE(n364),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][4] ),
	.D(n127),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][3]  (
	.SI(\REG_FILE[6][2] ),
	.SE(n426),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][3] ),
	.D(n126),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][2]  (
	.SI(\REG_FILE[6][1] ),
	.SE(n363),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][2] ),
	.D(n125),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][1]  (
	.SI(\REG_FILE[6][0] ),
	.SE(n425),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][1] ),
	.D(n124),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[6][0]  (
	.SI(\REG_FILE[5][7] ),
	.SE(n362),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[6][0] ),
	.D(n123),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][7]  (
	.SI(\REG_FILE[10][6] ),
	.SE(n318),
	.RN(RST),
	.Q(\REG_FILE[10][7] ),
	.D(n98),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][6]  (
	.SI(\REG_FILE[10][5] ),
	.SE(n380),
	.RN(RST),
	.Q(\REG_FILE[10][6] ),
	.D(n97),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][5]  (
	.SI(\REG_FILE[10][4] ),
	.SE(n317),
	.RN(RST),
	.Q(\REG_FILE[10][5] ),
	.D(n96),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][4]  (
	.SI(\REG_FILE[10][3] ),
	.SE(n379),
	.RN(RST),
	.Q(\REG_FILE[10][4] ),
	.D(n95),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][3]  (
	.SI(\REG_FILE[10][2] ),
	.SE(n316),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[10][3] ),
	.D(n94),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][2]  (
	.SI(\REG_FILE[10][1] ),
	.SE(n378),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[10][2] ),
	.D(n93),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][1]  (
	.SI(\REG_FILE[10][0] ),
	.SE(n300),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[10][1] ),
	.D(n92),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[10][0]  (
	.SI(\REG_FILE[9][7] ),
	.SE(n284),
	.RN(RST),
	.Q(\REG_FILE[10][0] ),
	.D(n91),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][7]  (
	.SI(\REG_FILE[14][6] ),
	.SE(n334),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[14][7] ),
	.D(n66),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][6]  (
	.SI(\REG_FILE[14][5] ),
	.SE(n396),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[14][6] ),
	.D(n65),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][5]  (
	.SI(\REG_FILE[14][4] ),
	.SE(n333),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[14][5] ),
	.D(n64),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][4]  (
	.SI(\REG_FILE[14][3] ),
	.SE(n395),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[14][4] ),
	.D(n63),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][3]  (
	.SI(\REG_FILE[14][2] ),
	.SE(n332),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[14][3] ),
	.D(n62),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][2]  (
	.SI(\REG_FILE[14][1] ),
	.SE(n394),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[14][2] ),
	.D(n61),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][1]  (
	.SI(\REG_FILE[14][0] ),
	.SE(n331),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[14][1] ),
	.D(n60),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[14][0]  (
	.SI(\REG_FILE[13][7] ),
	.SE(n393),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[14][0] ),
	.D(n59),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][7]  (
	.SI(\REG_FILE[4][6] ),
	.SE(n420),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][7] ),
	.D(n146),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][6]  (
	.SI(\REG_FILE[4][5] ),
	.SE(n357),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][6] ),
	.D(n145),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][5]  (
	.SI(\REG_FILE[4][4] ),
	.SE(n419),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][5] ),
	.D(n144),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][4]  (
	.SI(\REG_FILE[4][3] ),
	.SE(n356),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][4] ),
	.D(n143),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][3]  (
	.SI(\REG_FILE[4][2] ),
	.SE(n418),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][3] ),
	.D(n142),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][2]  (
	.SI(\REG_FILE[4][1] ),
	.SE(n355),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][2] ),
	.D(n141),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][1]  (
	.SI(\REG_FILE[4][0] ),
	.SE(n417),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][1] ),
	.D(n140),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[4][0]  (
	.SI(n472),
	.SE(n354),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[4][0] ),
	.D(n139),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][7]  (
	.SI(\REG_FILE[8][6] ),
	.SE(n315),
	.RN(RST),
	.Q(\REG_FILE[8][7] ),
	.D(n114),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][6]  (
	.SI(\REG_FILE[8][5] ),
	.SE(n304),
	.RN(RST),
	.Q(\REG_FILE[8][6] ),
	.D(n113),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][5]  (
	.SI(\REG_FILE[8][4] ),
	.SE(n288),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[8][5] ),
	.D(n112),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][4]  (
	.SI(test_si2),
	.SE(n289),
	.RN(RST),
	.Q(\REG_FILE[8][4] ),
	.D(n111),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][2]  (
	.SI(\REG_FILE[8][1] ),
	.SE(n371),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[8][2] ),
	.D(n109),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][1]  (
	.SI(\REG_FILE[8][0] ),
	.SE(n433),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[8][1] ),
	.D(n108),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[8][0]  (
	.SI(\REG_FILE[7][7] ),
	.SE(n370),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[8][0] ),
	.D(n107),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][7]  (
	.SI(\REG_FILE[12][6] ),
	.SE(n326),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][7] ),
	.D(n82),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][6]  (
	.SI(\REG_FILE[12][5] ),
	.SE(n388),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][6] ),
	.D(n81),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][5]  (
	.SI(\REG_FILE[12][4] ),
	.SE(n325),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][5] ),
	.D(n80),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][4]  (
	.SI(\REG_FILE[12][3] ),
	.SE(n387),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][4] ),
	.D(n79),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][3]  (
	.SI(\REG_FILE[12][2] ),
	.SE(n324),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][3] ),
	.D(n78),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][2]  (
	.SI(\REG_FILE[12][1] ),
	.SE(n386),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][2] ),
	.D(n77),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][1]  (
	.SI(\REG_FILE[12][0] ),
	.SE(n323),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[12][1] ),
	.D(n76),
	.CK(O_CLK1__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[12][0]  (
	.SI(\REG_FILE[11][7] ),
	.SE(n385),
	.RN(FE_OFN3_O_RST2),
	.Q(\REG_FILE[12][0] ),
	.D(n75),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[0]  (
	.SI(Rd_DATA_VLD),
	.SE(n339),
	.RN(FE_OFN3_O_RST2),
	.Q(Rd_DATA[0]),
	.D(n43),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][0]  (
	.SI(REG2[7]),
	.SE(n413),
	.RN(FE_OFN3_O_RST2),
	.Q(REG3[0]),
	.D(n147),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[2][1]  (
	.SI(REG2[0]),
	.SE(n412),
	.RN(FE_OFN3_O_RST2),
	.Q(REG2[1]),
	.D(n156),
	.CK(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[7]  (
	.SI(Rd_DATA[6]),
	.SE(n405),
	.RN(FE_OFN3_O_RST2),
	.Q(Rd_DATA[7]),
	.D(n50),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[6]  (
	.SI(Rd_DATA[5]),
	.SE(n342),
	.RN(FE_OFN3_O_RST2),
	.Q(Rd_DATA[6]),
	.D(n49),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[5]  (
	.SI(Rd_DATA[4]),
	.SE(n404),
	.RN(FE_OFN2_O_RST2),
	.Q(Rd_DATA[5]),
	.D(n48),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[4]  (
	.SI(Rd_DATA[3]),
	.SE(n341),
	.RN(FE_OFN3_O_RST2),
	.Q(Rd_DATA[4]),
	.D(n47),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[3]  (
	.SI(Rd_DATA[2]),
	.SE(n403),
	.RN(FE_OFN2_O_RST2),
	.Q(Rd_DATA[3]),
	.D(n46),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[2]  (
	.SI(Rd_DATA[1]),
	.SE(n340),
	.RN(FE_OFN2_O_RST2),
	.Q(Rd_DATA[2]),
	.D(n45),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Rd_DATA_reg[1]  (
	.SI(Rd_DATA[0]),
	.SE(n402),
	.RN(FE_OFN3_O_RST2),
	.Q(Rd_DATA[1]),
	.D(n44),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \REG_FILE_reg[3][5]  (
	.SN(RST),
	.SI(n474),
	.SE(n305),
	.Q(REG3[5]),
	.D(n152),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][2]  (
	.SI(n477),
	.SE(n414),
	.RN(FE_OFN3_O_RST2),
	.Q(n476),
	.D(n149),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][3]  (
	.SI(n476),
	.SE(n352),
	.RN(FE_OFN3_O_RST2),
	.Q(n475),
	.D(n150),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][4]  (
	.SI(n475),
	.SE(n415),
	.RN(FE_OFN3_O_RST2),
	.Q(n474),
	.D(n151),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \REG_FILE_reg[2][0]  (
	.SN(FE_OFN3_O_RST2),
	.SI(REG1[7]),
	.SE(n304),
	.Q(REG2[0]),
	.D(n155),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][7]  (
	.SI(n473),
	.SE(n416),
	.RN(RST),
	.Q(n472),
	.D(n154),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][6]  (
	.SI(REG3[5]),
	.SE(n353),
	.RN(FE_OFN3_O_RST2),
	.Q(n473),
	.D(n153),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[3][1]  (
	.SI(REG3[0]),
	.SE(n351),
	.RN(FE_OFN3_O_RST2),
	.Q(n477),
	.D(n148),
	.CK(O_CLK1__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][2]  (
	.SI(REG0[1]),
	.SE(n344),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[2]),
	.D(n173),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][0]  (
	.SI(test_si1),
	.SE(n343),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[0]),
	.D(n171),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][1]  (
	.SI(REG0[0]),
	.SE(n406),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[1]),
	.D(n172),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][5]  (
	.SI(REG0[4]),
	.SE(n408),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[5]),
	.D(n176),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][6]  (
	.SI(REG0[5]),
	.SE(n346),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[6]),
	.D(n177),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][7]  (
	.SI(REG0[6]),
	.SE(n409),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[7]),
	.D(n178),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[1][4]  (
	.SI(REG1[3]),
	.SE(n410),
	.RN(FE_OFN3_O_RST2),
	.Q(REG1[4]),
	.D(n167),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[1][5]  (
	.SI(REG1[4]),
	.SE(n348),
	.RN(FE_OFN3_O_RST2),
	.Q(REG1[5]),
	.D(n168),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[1][6]  (
	.SI(REG1[5]),
	.SE(n411),
	.RN(FE_OFN3_O_RST2),
	.Q(REG1[6]),
	.D(n169),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[1][7]  (
	.SI(REG1[6]),
	.SE(n349),
	.RN(FE_OFN3_O_RST2),
	.Q(REG1[7]),
	.D(n170),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][3]  (
	.SI(REG0[2]),
	.SE(n407),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[3]),
	.D(n174),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[0][4]  (
	.SI(REG0[3]),
	.SE(n345),
	.RN(FE_OFN3_O_RST2),
	.Q(REG0[4]),
	.D(n175),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[2][3]  (
	.SI(REG2[2]),
	.SE(n350),
	.RN(FE_OFN3_O_RST2),
	.Q(REG2[3]),
	.D(n158),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M Rd_DATA_VLD_reg (
	.SI(\REG_FILE[15][7] ),
	.SE(n401),
	.RN(FE_OFN3_O_RST2),
	.Q(Rd_DATA_VLD),
	.D(n42),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_FILE_reg[1][1]  (
	.SI(REG1[0]),
	.SE(n347),
	.RN(FE_OFN3_O_RST2),
	.Q(n275),
	.D(n164),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U61 (
	.Y(n281),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U285 (
	.Y(n282),
	.A(n299), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U286 (
	.Y(n283),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U287 (
	.Y(n284),
	.A(n377), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U288 (
	.Y(n285),
	.A(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U289 (
	.Y(n286),
	.A(n376), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U290 (
	.Y(n287),
	.A(n299), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U291 (
	.Y(n288),
	.A(n297), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U292 (
	.Y(n289),
	.A(n282), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U293 (
	.Y(REG3[1]),
	.A(n477), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U294 (
	.Y(REG3[7]),
	.A(n472), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U295 (
	.Y(REG3[3]),
	.A(n475), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U296 (
	.Y(REG3[2]),
	.A(n476), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U297 (
	.Y(REG3[4]),
	.A(n474), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U298 (
	.Y(n295),
	.A(n302), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U299 (
	.Y(n296),
	.A(n303), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U300 (
	.Y(n297),
	.A(n281), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U301 (
	.Y(n298),
	.A(n281), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U302 (
	.Y(n299),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U303 (
	.Y(n300),
	.A(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U304 (
	.Y(n306),
	.A(n282), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U305 (
	.Y(n301),
	.A(n306), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U306 (
	.Y(n309),
	.A(n283), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U307 (
	.Y(n302),
	.A(n309), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U308 (
	.Y(n308),
	.A(n297), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U309 (
	.Y(n303),
	.A(n308), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U310 (
	.Y(n304),
	.A(n283), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U311 (
	.Y(n305),
	.A(n298), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U312 (
	.Y(n307),
	.A(n298), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U316 (
	.Y(REG3[6]),
	.A(n473), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U317 (
	.Y(n314),
	.A(n286), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U318 (
	.Y(n315),
	.A(n284), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U319 (
	.Y(n316),
	.A(n378), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U320 (
	.Y(n317),
	.A(n379), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U321 (
	.Y(n318),
	.A(n380), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U322 (
	.Y(n319),
	.A(n381), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U323 (
	.Y(n320),
	.A(n382), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U324 (
	.Y(n321),
	.A(n383), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U325 (
	.Y(n322),
	.A(n384), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U326 (
	.Y(n323),
	.A(n385), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U327 (
	.Y(n324),
	.A(n386), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U328 (
	.Y(n325),
	.A(n387), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U329 (
	.Y(n326),
	.A(n388), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U330 (
	.Y(n327),
	.A(n389), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U331 (
	.Y(n328),
	.A(n390), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U332 (
	.Y(n329),
	.A(n391), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U333 (
	.Y(n330),
	.A(n392), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U334 (
	.Y(n331),
	.A(n393), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U335 (
	.Y(n332),
	.A(n394), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U336 (
	.Y(n333),
	.A(n395), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U337 (
	.Y(n334),
	.A(n396), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U338 (
	.Y(n335),
	.A(n397), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U339 (
	.Y(n336),
	.A(n398), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U340 (
	.Y(n337),
	.A(n399), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U341 (
	.Y(n338),
	.A(n400), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U342 (
	.Y(n339),
	.A(n401), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U343 (
	.Y(n340),
	.A(n402), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U344 (
	.Y(n341),
	.A(n403), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U345 (
	.Y(n342),
	.A(n404), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U346 (
	.Y(n343),
	.A(n405), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U347 (
	.Y(n344),
	.A(n406), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U348 (
	.Y(n345),
	.A(n407), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U349 (
	.Y(n346),
	.A(n408), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U350 (
	.Y(n347),
	.A(n409), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U351 (
	.Y(n348),
	.A(n410), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U352 (
	.Y(n349),
	.A(n411), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U353 (
	.Y(n350),
	.A(n412), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U354 (
	.Y(n351),
	.A(n413), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U355 (
	.Y(n352),
	.A(n414), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U356 (
	.Y(n353),
	.A(n415), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U357 (
	.Y(n354),
	.A(n416), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U358 (
	.Y(n355),
	.A(n417), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U359 (
	.Y(n356),
	.A(n418), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U360 (
	.Y(n357),
	.A(n419), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U361 (
	.Y(n358),
	.A(n420), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U362 (
	.Y(n359),
	.A(n421), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U363 (
	.Y(n360),
	.A(n422), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U364 (
	.Y(n361),
	.A(n423), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U365 (
	.Y(n362),
	.A(n424), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U366 (
	.Y(n363),
	.A(n425), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U367 (
	.Y(n364),
	.A(n426), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U368 (
	.Y(n365),
	.A(n427), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U369 (
	.Y(n366),
	.A(n428), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U370 (
	.Y(n367),
	.A(n429), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U371 (
	.Y(n368),
	.A(n430), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U372 (
	.Y(n369),
	.A(n431), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U373 (
	.Y(n370),
	.A(n432), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U374 (
	.Y(n371),
	.A(n433), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U379 (
	.Y(n376),
	.A(n287), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U380 (
	.Y(n377),
	.A(n285), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U381 (
	.Y(n378),
	.A(n300), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U382 (
	.Y(n379),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U383 (
	.Y(n380),
	.A(n317), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U384 (
	.Y(n381),
	.A(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U385 (
	.Y(n382),
	.A(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U386 (
	.Y(n383),
	.A(n320), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U387 (
	.Y(n384),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U388 (
	.Y(n385),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U389 (
	.Y(n386),
	.A(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U390 (
	.Y(n387),
	.A(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U391 (
	.Y(n388),
	.A(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U392 (
	.Y(n389),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U393 (
	.Y(n390),
	.A(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U394 (
	.Y(n391),
	.A(n328), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U395 (
	.Y(n392),
	.A(n329), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U396 (
	.Y(n393),
	.A(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U397 (
	.Y(n394),
	.A(n331), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U398 (
	.Y(n395),
	.A(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U399 (
	.Y(n396),
	.A(n333), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U400 (
	.Y(n397),
	.A(n334), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U401 (
	.Y(n398),
	.A(n335), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U402 (
	.Y(n399),
	.A(n336), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U403 (
	.Y(n400),
	.A(n337), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U404 (
	.Y(n401),
	.A(n338), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U405 (
	.Y(n402),
	.A(n339), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U406 (
	.Y(n403),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U407 (
	.Y(n404),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U408 (
	.Y(n405),
	.A(n342), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U409 (
	.Y(n406),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U410 (
	.Y(n407),
	.A(n344), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U411 (
	.Y(n408),
	.A(n345), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U412 (
	.Y(n409),
	.A(n346), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U413 (
	.Y(n410),
	.A(n347), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U414 (
	.Y(n411),
	.A(n348), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U415 (
	.Y(n412),
	.A(n349), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U416 (
	.Y(n413),
	.A(n350), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U417 (
	.Y(n414),
	.A(n351), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U418 (
	.Y(n415),
	.A(n352), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U419 (
	.Y(n416),
	.A(n353), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U420 (
	.Y(n417),
	.A(n354), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U421 (
	.Y(n418),
	.A(n355), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U422 (
	.Y(n419),
	.A(n356), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U423 (
	.Y(n420),
	.A(n357), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U424 (
	.Y(n421),
	.A(n358), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U425 (
	.Y(n422),
	.A(n359), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U426 (
	.Y(n423),
	.A(n360), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U427 (
	.Y(n424),
	.A(n361), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U428 (
	.Y(n425),
	.A(n362), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U429 (
	.Y(n426),
	.A(n363), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U430 (
	.Y(n427),
	.A(n364), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U431 (
	.Y(n428),
	.A(n365), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U432 (
	.Y(n429),
	.A(n366), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U433 (
	.Y(n430),
	.A(n367), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U434 (
	.Y(n431),
	.A(n368), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U435 (
	.Y(n432),
	.A(n369), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U436 (
	.Y(n433),
	.A(n370), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U438 (
	.Y(REG1[3]),
	.A(n434), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U439 (
	.Y(n436),
	.A(n466), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U440 (
	.Y(REG1[0]),
	.A(n436), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX1M \REG_FILE_reg[2][6]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(REG2[5]),
	.SE(n307),
	.RN(FE_OFN3_O_RST2),
	.Q(REG2[6]),
	.D(n161),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX1M \REG_FILE_reg[2][4]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(REG2[3]),
	.SE(n295),
	.RN(FE_OFN3_O_RST2),
	.Q(REG2[4]),
	.D(n159),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX1M \REG_FILE_reg[2][2]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(REG2[1]),
	.SE(n307),
	.RN(FE_OFN3_O_RST2),
	.Q(REG2[2]),
	.D(n157),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX1M \REG_FILE_reg[1][3]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(REG1[2]),
	.SE(n295),
	.RN(FE_OFN3_O_RST2),
	.QN(n434),
	.D(n166),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSRX1M \REG_FILE_reg[1][2]  (
	.SN(HTIE_LTIEHI_NET),
	.SI(REG1[1]),
	.SE(n296),
	.RN(FE_OFN3_O_RST2),
	.Q(REG1[2]),
	.D(n165),
	.CK(O_CLK1__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSX1M \REG_FILE_reg[2][7]  (
	.SN(FE_OFN3_O_RST2),
	.SI(REG2[6]),
	.SE(n289),
	.QN(n3),
	.D(n162),
	.CK(O_CLK1__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \REG_FILE_reg[8][3]  (
	.SI(\REG_FILE[8][2] ),
	.SE(n371),
	.RN(FE_OFN1_O_RST2),
	.Q(\REG_FILE[8][3] ),
	.D(n110),
	.CK(O_CLK1__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U6 (
	.Y(n2),
	.A(\REG_FILE[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX8M U437 (
	.Y(test_so1),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OUT_WD16_DATA_WD8_FUN_WD4_test_1 (
	A, 
	B, 
	ALU_FUN, 
	CLK, 
	RST, 
	ENABLE, 
	ALU_OUT, 
	OUT_VALID, 
	test_si, 
	test_se, 
	FE_OFN3_O_RST2, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input CLK;
   input RST;
   input ENABLE;
   output [15:0] ALU_OUT;
   output OUT_VALID;
   input test_si;
   input test_se;
   input FE_OFN3_O_RST2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_UNCONNECTED_0;
   wire n209;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N132;
   wire N133;
   wire N166;
   wire N168;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n186;
   wire n187;
   wire n188;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n210;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n56;

   // Module instantiations
   OAI2BB1X2M U11 (
	.Y(n61),
	.B0(n125),
	.A1N(n129),
	.A0N(n119), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U15 (
	.Y(n141),
	.B1(n195),
	.B0(n77),
	.A1N(n195),
	.A0N(ALU_OUT[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U16 (
	.Y(n140),
	.B1(n195),
	.B0(n63),
	.A1N(n195),
	.A0N(ALU_OUT[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U17 (
	.Y(n139),
	.B1(n46),
	.B0(ENABLE),
	.A1(n195),
	.A0(ALU_OUT[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n24),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U19 (
	.Y(n167),
	.B0(n164),
	.A1N(n166),
	.A0(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n176),
	.A(n167), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U21 (
	.Y(n26),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n170),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n169),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n168),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U25 (
	.Y(n88),
	.C1(n170),
	.C0(n90),
	.B1(n54),
	.B0(N129),
	.A1(n89),
	.A0(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U26 (
	.Y(n161),
	.B(B[6]),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U27 (
	.Y(n81),
	.C1(n169),
	.C0(n83),
	.B1(n54),
	.B0(N128),
	.A1(n82),
	.A0(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U28 (
	.Y(n95),
	.C1(n193),
	.C0(n97),
	.B1(n54),
	.B0(N130),
	.A1(n96),
	.A0(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U29 (
	.Y(n44),
	.B0(n155),
	.A2(n41),
	.A1(n42),
	.A0(n154), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U30 (
	.Y(n41),
	.C0(n40),
	.B0(n151),
	.A1(n172),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U31 (
	.Y(n109),
	.C1(n171),
	.C0(n111),
	.B1(n54),
	.B0(N132),
	.A1(n110),
	.A0(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U32 (
	.Y(n153),
	.C0(n150),
	.B0(n151),
	.A1(n173),
	.A0(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U33 (
	.Y(n151),
	.B(n156),
	.AN(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U34 (
	.Y(N168),
	.B0(n165),
	.A1(n149),
	.A0(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U35 (
	.Y(n102),
	.C1(n192),
	.C0(n104),
	.B1(n210),
	.B0(N131),
	.A1(n103),
	.A0(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U37 (
	.Y(n42),
	.B(A[2]),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U38 (
	.Y(n39),
	.B(A[0]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U39 (
	.Y(n154),
	.B(A[3]),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U42 (
	.Y(n68),
	.B(n129),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U43 (
	.Y(n69),
	.B(n76),
	.A(n119), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U44 (
	.Y(n123),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U45 (
	.Y(n119),
	.B(ALU_FUN[3]),
	.A(n206), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U46 (
	.Y(n124),
	.B(ALU_FUN[0]),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U47 (
	.Y(n76),
	.B(ALU_FUN[1]),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U49 (
	.Y(n186),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U50 (
	.Y(n164),
	.B(B[7]),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U54 (
	.Y(n199),
	.A(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U55 (
	.Y(n198),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U56 (
	.Y(n197),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U57 (
	.Y(n200),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U58 (
	.Y(n62),
	.B0(n125),
	.A1N(n124),
	.A0N(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U59 (
	.Y(n129),
	.B(n204),
	.A(n205), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U60 (
	.Y(n184),
	.A(n127), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U61 (
	.Y(n52),
	.B(n119),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U62 (
	.Y(n202),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U63 (
	.Y(n201),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U64 (
	.Y(n53),
	.B(n124),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U65 (
	.Y(n203),
	.A(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U68 (
	.Y(n55),
	.D(n206),
	.C(n76),
	.B(ALU_FUN[3]),
	.A(N168), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U69 (
	.Y(n173),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U70 (
	.Y(n107),
	.C1(n200),
	.C0(n27),
	.B1(n26),
	.B0(n197),
	.A1(n51),
	.A0(N114), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U71 (
	.Y(n114),
	.B1(n51),
	.B0(N115),
	.A1(n200),
	.A0(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U72 (
	.Y(n206),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U73 (
	.Y(n204),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U74 (
	.Y(n125),
	.C(n123),
	.B(ALU_FUN[3]),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U75 (
	.Y(n205),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U76 (
	.Y(n73),
	.C(n123),
	.B(n206),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U77 (
	.Y(n79),
	.C1(n200),
	.C0(A[2]),
	.B1(n188),
	.B0(n197),
	.A1(n51),
	.A0(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U78 (
	.Y(n86),
	.C1(n200),
	.C0(A[3]),
	.B1(n187),
	.B0(n197),
	.A1(n51),
	.A0(N111), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U79 (
	.Y(n93),
	.C1(n200),
	.C0(A[4]),
	.B1(n186),
	.B0(n197),
	.A1(n51),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U80 (
	.Y(n100),
	.C1(n200),
	.C0(A[5]),
	.B1(n24),
	.B0(n197),
	.A1(n51),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U81 (
	.Y(n127),
	.B0(ENABLE),
	.A1(n138),
	.A0(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U82 (
	.Y(n138),
	.B0(n197),
	.A1(n52),
	.A0(N107), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U83 (
	.Y(n196),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U85 (
	.Y(n51),
	.C(n204),
	.B(ALU_FUN[1]),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U86 (
	.Y(n175),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U87 (
	.Y(n60),
	.C(ALU_FUN[0]),
	.B(n76),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U88 (
	.Y(n72),
	.C(n129),
	.B(n206),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U89 (
	.Y(n131),
	.B(ENABLE),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U91 (
	.Y(n188),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U92 (
	.Y(n187),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U94 (
	.Y(n195),
	.A(ENABLE), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U99 (
	.Y(n57),
	.B(ALU_FUN[1]),
	.A(N166), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U100 (
	.Y(n74),
	.B0(n220),
	.A2(n75),
	.A1(ALU_FUN[0]),
	.A0(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U101 (
	.Y(n75),
	.C(n196),
	.B(ALU_FUN[2]),
	.A(n205), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U102 (
	.Y(n25),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U107 (
	.Y(n193),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U108 (
	.Y(n96),
	.C0(n69),
	.B1(n73),
	.B0(A[4]),
	.A1(n186),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U109 (
	.Y(n97),
	.C0(n68),
	.B1(n186),
	.B0(n73),
	.A1(n199),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U110 (
	.Y(n171),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U111 (
	.Y(n172),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U112 (
	.Y(n174),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U113 (
	.Y(n192),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U114 (
	.Y(n103),
	.C0(n69),
	.B1(n73),
	.B0(n25),
	.A1(n24),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U115 (
	.Y(n104),
	.C0(n68),
	.B1(n24),
	.B0(n73),
	.A1(n199),
	.A0(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U120 (
	.Y(n110),
	.C0(n69),
	.B1(n73),
	.B0(n27),
	.A1(n26),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U121 (
	.Y(n111),
	.C0(n68),
	.B1(n26),
	.B0(n73),
	.A1(n199),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U122 (
	.Y(n116),
	.C1(n191),
	.C0(n118),
	.B1(n54),
	.B0(N133),
	.A1(n117),
	.A0(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U123 (
	.Y(n191),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U124 (
	.Y(n117),
	.C0(n69),
	.B1(n73),
	.B0(A[7]),
	.A1(n175),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U125 (
	.Y(n118),
	.C0(n68),
	.B1(n175),
	.B0(n73),
	.A1(n199),
	.A0(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U126 (
	.Y(n66),
	.C1(n72),
	.C0(n190),
	.B1(n71),
	.B0(B[1]),
	.A1(n194),
	.A0(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U127 (
	.Y(n194),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U128 (
	.Y(n70),
	.C0(n200),
	.B1(n62),
	.B0(A[1]),
	.A1(n173),
	.A0(n202), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U129 (
	.Y(n71),
	.C0(n197),
	.B1(n173),
	.B0(n61),
	.A1(n202),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U130 (
	.Y(n27),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U132 (
	.Y(n190),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U134 (
	.Y(n49),
	.B1(n53),
	.B0(N90),
	.A1(n52),
	.A0(N99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U135 (
	.Y(n50),
	.C1(A[0]),
	.C0(n200),
	.B1(n190),
	.B0(n197),
	.A1(n51),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U136 (
	.Y(n63),
	.D(n67),
	.C(n66),
	.B(n65),
	.AN(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U137 (
	.Y(n64),
	.C1(n52),
	.C0(N100),
	.B1(n51),
	.B0(N109),
	.A1(n53),
	.A0(N91), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U138 (
	.Y(n67),
	.C1(n69),
	.C0(n173),
	.B1(n188),
	.B0(n60),
	.A1(n68),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U139 (
	.Y(n82),
	.C0(n69),
	.B1(n73),
	.B0(A[2]),
	.A1(n188),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U140 (
	.Y(n83),
	.C0(n68),
	.B1(n188),
	.B0(n73),
	.A1(n199),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4XLM U141 (
	.Y(n77),
	.D(n81),
	.C(n80),
	.B(n79),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U142 (
	.Y(n78),
	.B1(n53),
	.B0(N92),
	.A1(n52),
	.A0(N101), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U143 (
	.Y(n80),
	.B1(n203),
	.B0(A[3]),
	.A1(A[1]),
	.A0(n201), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U144 (
	.Y(n177),
	.A(n137), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U145 (
	.Y(n137),
	.C0(n184),
	.B1(n131),
	.B0(N123),
	.A1(n195),
	.A0(ALU_OUT[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U146 (
	.Y(n89),
	.C0(n69),
	.B1(n73),
	.B0(A[3]),
	.A1(n187),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U147 (
	.Y(n90),
	.C0(n68),
	.B1(n187),
	.B0(n73),
	.A1(n199),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n142),
	.B1(n195),
	.B0(n84),
	.A1N(n195),
	.A0N(ALU_OUT[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4XLM U149 (
	.Y(n84),
	.D(n88),
	.C(n87),
	.B(n86),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U150 (
	.Y(n85),
	.B1(n53),
	.B0(N93),
	.A1(n52),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U151 (
	.Y(n87),
	.B1(n203),
	.B0(A[4]),
	.A1(n201),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U152 (
	.Y(n178),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U153 (
	.Y(n136),
	.C0(n184),
	.B1(n131),
	.B0(N122),
	.A1(n195),
	.A0(ALU_OUT[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U156 (
	.Y(n143),
	.B1(n195),
	.B0(n91),
	.A1N(n195),
	.A0N(ALU_OUT[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4XLM U157 (
	.Y(n91),
	.D(n95),
	.C(n94),
	.B(n93),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U158 (
	.Y(n92),
	.B1(n53),
	.B0(N94),
	.A1(n52),
	.A0(N103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U159 (
	.Y(n94),
	.B1(n203),
	.B0(A[5]),
	.A1(n201),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U160 (
	.Y(n180),
	.A(n134), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U161 (
	.Y(n134),
	.C0(n184),
	.B1(n131),
	.B0(N120),
	.A1(n195),
	.A0(ALU_OUT[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U162 (
	.Y(n179),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U163 (
	.Y(n135),
	.C0(n184),
	.B1(n131),
	.B0(N121),
	.A1(n195),
	.A0(ALU_OUT[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U164 (
	.Y(n144),
	.B1(n195),
	.B0(n98),
	.A1N(n195),
	.A0N(ALU_OUT[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4XLM U165 (
	.Y(n98),
	.D(n102),
	.C(n101),
	.B(n100),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U166 (
	.Y(n99),
	.B1(n53),
	.B0(N95),
	.A1(n52),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U167 (
	.Y(n101),
	.B1(n203),
	.B0(n27),
	.A1(n201),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U168 (
	.Y(n182),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U169 (
	.Y(n132),
	.C0(n184),
	.B1(n131),
	.B0(N118),
	.A1(n195),
	.A0(ALU_OUT[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U170 (
	.Y(n181),
	.A(n133), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U171 (
	.Y(n133),
	.C0(n184),
	.B1(n131),
	.B0(N119),
	.A1(n195),
	.A0(ALU_OUT[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U172 (
	.Y(n54),
	.C(n120),
	.B(ALU_FUN[1]),
	.A(n119), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U173 (
	.Y(n120),
	.B0(ALU_FUN[2]),
	.A1(n122),
	.A0(n121), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U174 (
	.Y(n122),
	.D(B[4]),
	.C(B[5]),
	.B(B[6]),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U175 (
	.Y(n121),
	.D(B[0]),
	.C(B[1]),
	.B(B[2]),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U176 (
	.Y(n147),
	.C0(n128),
	.B0(n127),
	.A1(n195),
	.A0(n126), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U177 (
	.Y(n128),
	.B(n195),
	.A(ALU_OUT[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U178 (
	.Y(n126),
	.C1(n51),
	.C0(N116),
	.B1(n201),
	.B0(A[7]),
	.A1(n53),
	.A0(N98), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U179 (
	.Y(n145),
	.B1(n195),
	.B0(n105),
	.A1N(n195),
	.A0N(ALU_OUT[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4XLM U180 (
	.Y(n105),
	.D(n109),
	.C(n108),
	.B(n107),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U181 (
	.Y(n106),
	.B1(n53),
	.B0(N96),
	.A1(n52),
	.A0(N105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U182 (
	.Y(n108),
	.B1(n203),
	.B0(A[7]),
	.A1(n201),
	.A0(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U183 (
	.Y(n146),
	.B1(n195),
	.B0(n112),
	.A1N(n195),
	.A0N(ALU_OUT[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U184 (
	.Y(n112),
	.D(n116),
	.C(n115),
	.B(n114),
	.A(n113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U185 (
	.Y(n113),
	.B1(n53),
	.B0(N97),
	.A1(n52),
	.A0(N106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U186 (
	.Y(n115),
	.B1(n175),
	.B0(n197),
	.A1(n201),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U187 (
	.Y(n183),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U188 (
	.Y(n130),
	.C0(n184),
	.B1(n131),
	.B0(N117),
	.A1(n195),
	.A0(ALU_OUT[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U189 (
	.Y(n47),
	.C1(n173),
	.C0(n60),
	.B1(n59),
	.B0(B[0]),
	.A1(n168),
	.A0(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U190 (
	.Y(n58),
	.C0(n200),
	.B1(n62),
	.B0(A[0]),
	.A1(n190),
	.A0(n202), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U191 (
	.Y(n59),
	.C0(n197),
	.B1(n190),
	.B0(n61),
	.A1(n202),
	.A0(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U192 (
	.Y(n148),
	.B(n195),
	.AN(n247), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1XLM U193 (
	.Y(n65),
	.B0(n74),
	.A1N(n54),
	.A0N(N127), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U194 (
	.Y(n157),
	.B(A[4]),
	.AN(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U195 (
	.Y(n43),
	.B(B[4]),
	.AN(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U196 (
	.Y(n159),
	.B(n43),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U197 (
	.Y(n156),
	.B(n169),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U198 (
	.Y(n40),
	.B0(B[1]),
	.A1(n173),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U199 (
	.Y(n155),
	.B(n170),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U200 (
	.Y(n162),
	.B(B[5]),
	.AN(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U201 (
	.Y(n45),
	.C0(n162),
	.B0(n43),
	.A1(n44),
	.A0(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U202 (
	.Y(n158),
	.B(n25),
	.AN(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U203 (
	.Y(n149),
	.B1(n26),
	.B0(B[6]),
	.A2(n161),
	.A1(n158),
	.A0(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U204 (
	.Y(n165),
	.B(n175),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U205 (
	.Y(n152),
	.B(n168),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U206 (
	.Y(n150),
	.B0(B[1]),
	.A1(n173),
	.A0(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U207 (
	.Y(n160),
	.B0(n154),
	.A2(n155),
	.A1(n156),
	.A0(n174), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X1M U208 (
	.Y(n163),
	.C0(n157),
	.B0(n158),
	.A1N(n160),
	.A0(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U209 (
	.Y(n166),
	.B1(n171),
	.B0(n27),
	.A2(n161),
	.A1(n162),
	.A0(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U210 (
	.Y(N166),
	.B(n176),
	.A(N168), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(n218),
	.RN(RST),
	.Q(ALU_OUT[7]),
	.D(n146),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(n221),
	.RN(RST),
	.Q(ALU_OUT[6]),
	.D(n145),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(n223),
	.RN(RST),
	.Q(ALU_OUT[5]),
	.D(n144),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(n217),
	.RN(RST),
	.Q(ALU_OUT[4]),
	.D(n143),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(n233),
	.RN(RST),
	.Q(ALU_OUT[3]),
	.D(n142),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(n222),
	.RN(FE_OFN3_O_RST2),
	.Q(ALU_OUT[1]),
	.D(n140),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(n219),
	.RN(RST),
	.Q(ALU_OUT[15]),
	.D(n177),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(n234),
	.RN(RST),
	.Q(ALU_OUT[14]),
	.D(n178),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(n223),
	.RN(RST),
	.Q(ALU_OUT[13]),
	.D(n179),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(n221),
	.RN(RST),
	.Q(ALU_OUT[12]),
	.D(n180),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(n218),
	.RN(RST),
	.Q(ALU_OUT[11]),
	.D(n181),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(n230),
	.RN(RST),
	.Q(ALU_OUT[10]),
	.D(n182),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(n222),
	.RN(RST),
	.Q(ALU_OUT[9]),
	.D(n183),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(n232),
	.RN(RST),
	.Q(ALU_OUT[8]),
	.D(n147),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M OUT_VALID_reg (
	.SI(ALU_OUT[15]),
	.SE(n219),
	.RN(FE_OFN3_O_RST2),
	.Q(n209),
	.D(n148),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(n216),
	.RN(RST),
	.Q(ALU_OUT[2]),
	.D(n141),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[0]  (
	.SI(test_si),
	.SE(n217),
	.RN(FE_OFN3_O_RST2),
	.Q(ALU_OUT[0]),
	.D(n139),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U36 (
	.Y(n210),
	.A(n244), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U214 (
	.Y(n215),
	.A(n229), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U215 (
	.Y(n216),
	.A(n232), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U216 (
	.Y(n217),
	.A(n230), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U217 (
	.Y(n218),
	.A(n233), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U218 (
	.Y(n219),
	.A(n234), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U219 (
	.Y(n220),
	.A(n245), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U220 (
	.Y(n221),
	.A(n229), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U221 (
	.Y(n222),
	.A(n231), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U222 (
	.Y(n223),
	.A(n231), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U226 (
	.Y(n227),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U227 (
	.Y(n228),
	.A(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U228 (
	.Y(n229),
	.A(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U229 (
	.Y(n230),
	.A(n215), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U230 (
	.Y(n231),
	.A(n228), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U231 (
	.Y(n232),
	.A(n215), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U232 (
	.Y(n233),
	.A(n228), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U233 (
	.Y(n234),
	.A(n216), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U234 (
	.Y(n235),
	.C(n241),
	.B(n49),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U235 (
	.Y(n46),
	.B(n236),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U236 (
	.Y(n236),
	.A(n235), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U241 (
	.Y(n241),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U242 (
	.Y(n242),
	.C0(n246),
	.B0(n245),
	.A1(n244),
	.A0(n243), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U243 (
	.Y(n48),
	.A(n242), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U244 (
	.Y(n243),
	.A(N126), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U245 (
	.Y(n244),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U246 (
	.Y(n245),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U247 (
	.Y(n246),
	.D(ALU_FUN[0]),
	.C(ALU_FUN[2]),
	.B(n196),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M U248 (
	.Y(n247),
	.A(OUT_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW_div_uns_0 div_29 (
	.a({ A[7],
		A[6],
		n25,
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.b({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		n169,
		B[1],
		B[0] }),
	.quotient({ N133,
		N132,
		N131,
		N130,
		N129,
		N128,
		N127,
		N126 }),
	.n169(n169),
	.n170(n170),
	.n194(n194),
	.n187(n187),
	.n191(n191),
	.n171(n171),
	.n192(n192),
	.n193(n193),
	.n173(n173),
	.n168(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW01_sub_0 sub_21 (
	.A({ 1'b0,
		A[7],
		n27,
		n25,
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.DIFF({ N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101,
		N100,
		N99 }),
	.n170(n170),
	.n194(n194),
	.n191(n191),
	.n171(n171),
	.n192(n192),
	.n193(n193),
	.n168(n168),
	.n169(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW01_add_0 add_18 (
	.A({ 1'b0,
		A[7],
		A[6],
		n25,
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.SUM({ N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92,
		N91,
		N90 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW02_mult_0 mult_24 (
	.A({ A[7],
		n27,
		n25,
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.TC(1'b0),
	.PRODUCT({ N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109,
		N108 }),
	.n169(n169),
	.n238(FE_UNCONNECTED_0),
	.n170(n170),
	.n194(n194),
	.n186(n186),
	.n187(n187),
	.n191(n191),
	.n171(n171),
	.n192(n192),
	.n193(n193),
	.n175(n175),
	.n173(n173),
	.n190(n190),
	.n188(n188),
	.n168(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U249 (
	.Y(n56),
	.A(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX8M U250 (
	.Y(OUT_VALID),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n169, 
	n170, 
	n194, 
	n187, 
	n191, 
	n171, 
	n192, 
	n193, 
	n173, 
	n168, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n169;
   input n170;
   input n194;
   input n187;
   input n191;
   input n171;
   input n192;
   input n193;
   input n173;
   input n168;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n25;
   wire n28;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[1][4] ;
   wire \u_div/CryTmp[1][5] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][4] ;
   wire \u_div/CryTmp[2][5] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[3][4] ;
   wire \u_div/CryTmp[3][5] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[4][4] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[6][2] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n6;
   wire n8;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n22;
   wire n23;
   wire n24;
   wire n34;
   wire n35;
   wire n38;
   wire n39;
   wire n41;
   wire n42;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n59;
   wire n61;

   // Module instantiations
   ADDFX2M \u_div/u_fa_PartRem_0_1_1  (
	.S(\u_div/SumTmp[1][1] ),
	.CO(\u_div/CryTmp[1][2] ),
	.CI(\u_div/PartRem[2][1] ),
	.B(n194),
	.A(\u_div/CryTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_1  (
	.S(\u_div/SumTmp[3][1] ),
	.CO(\u_div/CryTmp[3][2] ),
	.CI(\u_div/CryTmp[3][1] ),
	.B(n194),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_1  (
	.S(\u_div/SumTmp[4][1] ),
	.CO(\u_div/CryTmp[4][2] ),
	.CI(\u_div/CryTmp[4][1] ),
	.B(n194),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_3  (
	.S(\u_div/SumTmp[4][3] ),
	.CO(\u_div/CryTmp[4][4] ),
	.CI(\u_div/CryTmp[4][3] ),
	.B(n170),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/PartRem[1][1] ),
	.B(n194),
	.A(\u_div/CryTmp[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(n169),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(n170),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(n171),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_2  (
	.S(\u_div/SumTmp[3][2] ),
	.CO(\u_div/CryTmp[3][3] ),
	.CI(\u_div/CryTmp[3][2] ),
	.B(n169),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_2  (
	.S(\u_div/SumTmp[4][2] ),
	.CO(\u_div/CryTmp[4][3] ),
	.CI(\u_div/CryTmp[4][2] ),
	.B(n169),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_3  (
	.S(\u_div/SumTmp[3][3] ),
	.CO(\u_div/CryTmp[3][4] ),
	.CI(\u_div/CryTmp[3][3] ),
	.B(n170),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_6_1  (
	.S(\u_div/SumTmp[6][1] ),
	.CO(\u_div/CryTmp[6][2] ),
	.CI(\u_div/CryTmp[6][1] ),
	.B(n194),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_2  (
	.S(\u_div/SumTmp[1][2] ),
	.CO(\u_div/CryTmp[1][3] ),
	.CI(\u_div/CryTmp[1][2] ),
	.B(n169),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(n191),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_6  (
	.S(\u_div/SumTmp[1][6] ),
	.CO(\u_div/CryTmp[1][7] ),
	.CI(\u_div/CryTmp[1][6] ),
	.B(n171),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_3  (
	.S(\u_div/SumTmp[2][3] ),
	.CO(\u_div/CryTmp[2][4] ),
	.CI(\u_div/CryTmp[2][3] ),
	.B(n170),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_2  (
	.S(\u_div/SumTmp[2][2] ),
	.CO(\u_div/CryTmp[2][3] ),
	.CI(\u_div/CryTmp[2][2] ),
	.B(n169),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_1  (
	.S(\u_div/SumTmp[2][1] ),
	.CO(\u_div/CryTmp[2][2] ),
	.CI(\u_div/PartRem[3][1] ),
	.B(n194),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_5  (
	.S(\u_div/SumTmp[2][5] ),
	.CO(\u_div/CryTmp[2][6] ),
	.CI(\u_div/CryTmp[2][5] ),
	.B(n192),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_5  (
	.S(\u_div/SumTmp[1][5] ),
	.CO(\u_div/CryTmp[1][6] ),
	.CI(\u_div/CryTmp[1][5] ),
	.B(n192),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(n192),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_4  (
	.S(\u_div/SumTmp[2][4] ),
	.CO(\u_div/CryTmp[2][5] ),
	.CI(\u_div/CryTmp[2][4] ),
	.B(n193),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_4  (
	.S(\u_div/SumTmp[3][4] ),
	.CO(\u_div/CryTmp[3][5] ),
	.CI(\u_div/CryTmp[3][4] ),
	.B(n193),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_4  (
	.S(\u_div/SumTmp[1][4] ),
	.CO(\u_div/CryTmp[1][5] ),
	.CI(\u_div/CryTmp[1][4] ),
	.B(n193),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(n193),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_2  (
	.S(\u_div/SumTmp[5][2] ),
	.CO(\u_div/CryTmp[5][3] ),
	.CI(\u_div/CryTmp[5][2] ),
	.B(n169),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_1  (
	.S(\u_div/SumTmp[5][1] ),
	.CO(\u_div/CryTmp[5][2] ),
	.CI(\u_div/CryTmp[5][1] ),
	.B(n194),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(\u_div/PartRem[6][1] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][0] ),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U2 (
	.Y(\u_div/PartRem[5][1] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][0] ),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U4 (
	.Y(n24),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U7 (
	.Y(n11),
	.B(n10),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(n168),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(quotient[2]),
	.B(n24),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U11 (
	.Y(\u_div/PartRem[3][2] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][1] ),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U15 (
	.Y(\u_div/PartRem[6][2] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][1] ),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U16 (
	.Y(\u_div/PartRem[2][4] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U17 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][6] ),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U18 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U19 (
	.Y(n1),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U20 (
	.Y(quotient[1]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U22 (
	.Y(quotient[4]),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U23 (
	.Y(n28),
	.B(n191),
	.A(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U25 (
	.Y(\u_div/PartRem[3][3] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U30 (
	.Y(n6),
	.B(n24),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U31 (
	.Y(n23),
	.B(n6),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U33 (
	.Y(quotient[7]),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U34 (
	.Y(n10),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U35 (
	.Y(n25),
	.B(n8),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U36 (
	.Y(n22),
	.B(n170),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U37 (
	.Y(n8),
	.C(n194),
	.B(n169),
	.A(\u_div/CryTmp[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U38 (
	.Y(quotient[6]),
	.B(n13),
	.A(\u_div/CryTmp[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U39 (
	.Y(n12),
	.B(n25),
	.A(\u_div/SumTmp[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U40 (
	.Y(\u_div/PartRem[7][1] ),
	.B(n12),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U41 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][0] ),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U43 (
	.Y(n13),
	.B(b[2]),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U44 (
	.Y(\u_div/PartRem[4][2] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][1] ),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U45 (
	.Y(\u_div/PartRem[4][3] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][2] ),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U46 (
	.Y(\u_div/PartRem[3][4] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U47 (
	.Y(\u_div/SumTmp[5][0] ),
	.B(a[5]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U48 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U49 (
	.Y(\u_div/SumTmp[4][0] ),
	.B(a[4]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U51 (
	.Y(\u_div/SumTmp[6][0] ),
	.B(a[6]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U52 (
	.Y(\u_div/CryTmp[5][1] ),
	.B(n168),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U53 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(n168),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U54 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n168),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U55 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(a[1]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U57 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(n168),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U60 (
	.Y(\u_div/PartRem[5][2] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][1] ),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U61 (
	.Y(\u_div/CryTmp[4][1] ),
	.B(n168),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U62 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(b[0]),
	.AN(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U66 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][5] ),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U67 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][4] ),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U68 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][3] ),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U70 (
	.Y(\u_div/PartRem[2][6] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U71 (
	.Y(\u_div/PartRem[2][5] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U72 (
	.Y(\u_div/PartRem[3][5] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U73 (
	.Y(\u_div/PartRem[4][4] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U74 (
	.Y(\u_div/PartRem[5][3] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U28 (
	.Y(n48),
	.B(n34),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U29 (
	.Y(n34),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n35),
	.B(\u_div/CryTmp[4][4] ),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U65 (
	.Y(n38),
	.A(\u_div/CryTmp[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U69 (
	.Y(n39),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U75 (
	.Y(\u_div/PartRem[3][1] ),
	.S0(n59),
	.B(n187),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U77 (
	.Y(n41),
	.A(\u_div/SumTmp[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U78 (
	.Y(n42),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][0] ),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U79 (
	.Y(\u_div/PartRem[2][1] ),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U82 (
	.Y(n45),
	.B(n24),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U83 (
	.Y(n59),
	.B(n46),
	.A(\u_div/CryTmp[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U84 (
	.Y(n46),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U85 (
	.Y(n47),
	.B(\u_div/PartRem[2][3] ),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U86 (
	.Y(\u_div/SumTmp[1][3] ),
	.B(n39),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U87 (
	.Y(n49),
	.B(n170),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U88 (
	.Y(n50),
	.B(n170),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U89 (
	.Y(\u_div/CryTmp[1][4] ),
	.C(n48),
	.B(n49),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U90 (
	.Y(n51),
	.B(n22),
	.A(\u_div/CryTmp[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U91 (
	.Y(quotient[5]),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U92 (
	.Y(n52),
	.S0(quotient[1]),
	.B(n53),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U93 (
	.Y(\u_div/PartRem[1][3] ),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U94 (
	.Y(n53),
	.A(\u_div/SumTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U95 (
	.Y(n54),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][1] ),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U96 (
	.Y(\u_div/PartRem[2][2] ),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U97 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(n56),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U98 (
	.Y(n55),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U99 (
	.Y(n56),
	.A(\u_div/SumTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U102 (
	.Y(quotient[3]),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U103 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(n1),
	.B(n173),
	.A(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U105 (
	.Y(n61),
	.B(a[1]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n170, 
	n194, 
	n191, 
	n171, 
	n192, 
	n193, 
	n168, 
	n169, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n170;
   input n194;
   input n191;
   input n171;
   input n192;
   input n193;
   input n168;
   input n169;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n169),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n170),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n194),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n171),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n192),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n193),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n191),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(carry[1]),
	.B(n168),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U11 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U2 (
	.Y(SUM[0]),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n169, 
	n238, 
	n170, 
	n194, 
	n186, 
	n187, 
	n191, 
	n171, 
	n192, 
	n193, 
	n175, 
	n173, 
	n190, 
	n188, 
	n168, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n169;
   input n238;
   input n170;
   input n194;
   input n186;
   input n187;
   input n191;
   input n171;
   input n192;
   input n193;
   input n175;
   input n173;
   input n190;
   input n188;
   input n168;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n18;
   wire n19;

   // Module instantiations
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n9),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n7),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n4),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n8),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n6),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n5),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n3),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U10 (
	.Y(\ab[0][4] ),
	.B(n190),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U11 (
	.Y(\ab[0][7] ),
	.B(n190),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(\ab[0][5] ),
	.B(n190),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U13 (
	.Y(\ab[0][6] ),
	.B(n190),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U14 (
	.Y(\ab[0][1] ),
	.B(n190),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(\ab[1][6] ),
	.B(n173),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(\ab[1][4] ),
	.B(n173),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(\ab[1][5] ),
	.B(n173),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(\ab[1][1] ),
	.B(n173),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(\ab[7][7] ),
	.B(n191),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U20 (
	.Y(PRODUCT[1]),
	.B(\ab[0][1] ),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(\ab[0][3] ),
	.B(n190),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(\ab[1][3] ),
	.B(n173),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(\ab[1][2] ),
	.B(n173),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(\ab[0][2] ),
	.B(n190),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U25 (
	.Y(\ab[1][0] ),
	.B(n173),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U27 (
	.Y(n19),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U33 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U34 (
	.Y(n11),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U35 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U36 (
	.Y(n12),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U37 (
	.Y(n13),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U39 (
	.Y(\SUMB[1][2] ),
	.B(\ab[0][3] ),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U43 (
	.Y(n14),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U44 (
	.Y(\SUMB[1][5] ),
	.B(\ab[0][6] ),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U45 (
	.Y(\SUMB[1][6] ),
	.B(\ab[0][7] ),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U46 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U49 (
	.Y(n18),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U50 (
	.Y(n16),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(\A1[6] ),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U52 (
	.Y(\SUMB[1][3] ),
	.B(\ab[0][4] ),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U53 (
	.Y(\SUMB[1][4] ),
	.B(\ab[0][5] ),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U59 (
	.Y(\SUMB[1][1] ),
	.B(\ab[0][2] ),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[7][6] ),
	.B(n171),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[7][5] ),
	.B(n192),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[7][4] ),
	.B(n193),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[7][3] ),
	.B(n170),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[7][2] ),
	.B(n169),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[7][1] ),
	.B(n194),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[7][0] ),
	.B(n168),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][7] ),
	.B(n18),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[6][6] ),
	.B(n18),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[6][5] ),
	.B(n18),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[6][4] ),
	.B(n18),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[6][3] ),
	.B(n18),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[6][2] ),
	.B(n18),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[6][1] ),
	.B(n18),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[6][0] ),
	.B(n18),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][7] ),
	.B(n19),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[5][6] ),
	.B(n19),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[5][5] ),
	.B(n19),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[5][4] ),
	.B(n19),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[5][3] ),
	.B(n19),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[5][2] ),
	.B(n19),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[5][1] ),
	.B(n19),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[5][0] ),
	.B(n19),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][7] ),
	.B(n186),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[4][6] ),
	.B(n186),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[4][5] ),
	.B(n186),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[4][4] ),
	.B(n186),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[4][3] ),
	.B(n186),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[4][2] ),
	.B(n186),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[4][1] ),
	.B(n186),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[4][0] ),
	.B(n186),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][7] ),
	.B(n187),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[3][6] ),
	.B(n187),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[3][5] ),
	.B(n187),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[3][4] ),
	.B(n187),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[3][3] ),
	.B(n187),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[3][2] ),
	.B(n187),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[3][1] ),
	.B(n187),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[3][0] ),
	.B(n187),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][7] ),
	.B(n188),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[2][6] ),
	.B(n188),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[2][5] ),
	.B(n188),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[2][4] ),
	.B(n188),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[2][3] ),
	.B(n188),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[2][2] ),
	.B(n188),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[2][1] ),
	.B(n188),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[2][0] ),
	.B(n188),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][7] ),
	.B(n173),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(PRODUCT[0]),
	.B(n190),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n12,
		n11,
		n16,
		n15,
		n13,
		n14,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OUT_WD16_DATA_WD8_FUN_WD4_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;

   // Module instantiations
   OAI21BX1M U2 (
	.Y(n17),
	.B0N(n21),
	.A1(n20),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U3 (
	.Y(n24),
	.B0(n10),
	.A1N(n11),
	.A0N(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1XLM U4 (
	.Y(n16),
	.B0(n18),
	.A1N(A[12]),
	.A0N(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(n19),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n14),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(n11),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U8 (
	.Y(n23),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n13),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n7),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(SUM[13]),
	.B(n16),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(SUM[6]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(SUM[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U14 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U15 (
	.Y(SUM[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U16 (
	.Y(SUM[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U17 (
	.Y(SUM[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U18 (
	.Y(SUM[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U19 (
	.Y(SUM[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U20 (
	.Y(SUM[9]),
	.B(n9),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U21 (
	.Y(n9),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(SUM[8]),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U23 (
	.Y(n12),
	.B(n15),
	.AN(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U24 (
	.Y(n18),
	.B0(B[12]),
	.A1(n17),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U25 (
	.Y(SUM[12]),
	.C(n17),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U26 (
	.Y(SUM[11]),
	.B(n22),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U27 (
	.Y(n22),
	.B(n19),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U28 (
	.Y(n21),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U29 (
	.Y(n20),
	.B0(n25),
	.A1(n24),
	.A0(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(SUM[10]),
	.B(n24),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U31 (
	.Y(n10),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U32 (
	.Y(n8),
	.B0(n15),
	.A1(n14),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U33 (
	.Y(n15),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U34 (
	.Y(n26),
	.B(n25),
	.AN(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n25),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_GATE (
	CLK_EN, 
	CLK, 
	GATED_CLK, 
	VDD, 
	VSS);
   input CLK_EN;
   input CLK;
   output GATED_CLK;
   inout VDD;
   inout VSS;

   // Module instantiations
   TLATNCAX12M U0_TLATNCAX12M (
	.ECK(GATED_CLK),
	.E(CLK_EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_TOP (
	RST_N, 
	UART_CLK, 
	REF_CLK, 
	UART_RX_IN, 
	SI, 
	SE, 
	test_mode, 
	scan_clk, 
	scan_rst, 
	SO, 
	UART_TX_O, 
	parity_error, 
	framing_error, 
	VDD, 
	VSS);
   input RST_N;
   input UART_CLK;
   input REF_CLK;
   input UART_RX_IN;
   input [3:0] SI;
   input SE;
   input test_mode;
   input scan_clk;
   input scan_rst;
   output [3:0] SO;
   output UART_TX_O;
   output parity_error;
   output framing_error;
   inout VDD;
   inout VSS;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L14_N0;
   wire scan_clk__L13_N0;
   wire scan_clk__L12_N1;
   wire scan_clk__L12_N0;
   wire scan_clk__L11_N1;
   wire scan_clk__L11_N0;
   wire scan_clk__L10_N1;
   wire scan_clk__L10_N0;
   wire scan_clk__L9_N1;
   wire scan_clk__L9_N0;
   wire scan_clk__L8_N1;
   wire scan_clk__L8_N0;
   wire scan_clk__L7_N1;
   wire scan_clk__L7_N0;
   wire scan_clk__L6_N1;
   wire scan_clk__L6_N0;
   wire scan_clk__L5_N1;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N1;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire O_CLK1__L5_N7;
   wire O_CLK1__L5_N6;
   wire O_CLK1__L5_N5;
   wire O_CLK1__L5_N4;
   wire O_CLK1__L5_N3;
   wire O_CLK1__L5_N2;
   wire O_CLK1__L5_N1;
   wire O_CLK1__L5_N0;
   wire O_CLK1__L4_N3;
   wire O_CLK1__L4_N2;
   wire O_CLK1__L4_N1;
   wire O_CLK1__L4_N0;
   wire O_CLK1__L3_N1;
   wire O_CLK1__L3_N0;
   wire O_CLK1__L2_N0;
   wire O_CLK1__L1_N0;
   wire ALU_CLK__L3_N0;
   wire ALU_CLK__L2_N0;
   wire ALU_CLK__L1_N0;
   wire O_CLK2__L13_N0;
   wire O_CLK2__L12_N0;
   wire O_CLK2__L11_N0;
   wire O_CLK2__L10_N0;
   wire O_CLK2__L9_N0;
   wire O_CLK2__L8_N0;
   wire O_CLK2__L7_N1;
   wire O_CLK2__L7_N0;
   wire O_CLK2__L6_N1;
   wire O_CLK2__L6_N0;
   wire O_CLK2__L5_N0;
   wire O_CLK2__L4_N0;
   wire O_CLK2__L3_N0;
   wire O_CLK2__L2_N0;
   wire O_CLK2__L1_N0;
   wire O_CLK3__L3_N3;
   wire O_CLK3__L3_N2;
   wire O_CLK3__L3_N1;
   wire O_CLK3__L3_N0;
   wire O_CLK3__L2_N0;
   wire O_CLK3__L1_N0;
   wire O_CLK4__L3_N1;
   wire O_CLK4__L3_N0;
   wire O_CLK4__L2_N0;
   wire O_CLK4__L1_N0;
   wire FE_OFN3_O_RST2;
   wire FE_OFN2_O_RST2;
   wire FE_OFN0_O_RST2;
   wire O_CLK1;
   wire O_CLK2;
   wire TX_CLK;
   wire O_CLK3;
   wire RX_CLK;
   wire O_CLK4;
   wire O_RST1;
   wire SYNC_RST1;
   wire O_RST2;
   wire SYNC_RST2;
   wire O_RST3;
   wire RX_VLD;
   wire RX_VLD_SYNC;
   wire WR_INC;
   wire RD_INC;
   wire FIFO_FULL;
   wire F_EMPTY;
   wire BUSY;
   wire ALU_OUT_VLD;
   wire RD_D_VLD;
   wire ALU_EN;
   wire GATE_EN;
   wire WrEn;
   wire RdEn;
   wire ALU_CLK;
   wire _1_net_;
   wire n1;
   wire n2;
   wire n4;
   wire n5;
   wire n13;
   wire n14;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n23;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire [7:0] RX_OUT_P;
   wire [7:0] RX_OUT_SYNC;
   wire [7:0] WR_DATA;
   wire [7:0] RD_DATA;
   wire [7:0] div_ratio;
   wire [7:0] UART_CONFIG;
   wire [3:0] Pre_div;
   wire [15:0] ALU_OUT;
   wire [7:0] Rd_D;
   wire [3:0] ALU_FUN;
   wire [3:0] Address;
   wire [7:0] Wr_D;
   wire [7:0] Op_A;
   wire [7:0] Op_B;

   assign SO[0] = ALU_OUT_VLD ;

   // Module instantiations
   CLKINVX16M REF_CLK__L2_I0 (
	.Y(REF_CLK__L2_N0),
	.A(REF_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M REF_CLK__L1_I0 (
	.Y(REF_CLK__L1_N0),
	.A(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M UART_CLK__L2_I0 (
	.Y(UART_CLK__L2_N0),
	.A(UART_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_CLK__L1_I0 (
	.Y(UART_CLK__L1_N0),
	.A(UART_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk__L14_I0 (
	.Y(scan_clk__L14_N0),
	.A(scan_clk__L13_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L13_I0 (
	.Y(scan_clk__L13_N0),
	.A(scan_clk__L12_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk__L12_I1 (
	.Y(scan_clk__L12_N1),
	.A(scan_clk__L11_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX24M scan_clk__L12_I0 (
	.Y(scan_clk__L12_N0),
	.A(scan_clk__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L11_I1 (
	.Y(scan_clk__L11_N1),
	.A(scan_clk__L10_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L11_I0 (
	.Y(scan_clk__L11_N0),
	.A(scan_clk__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L10_I1 (
	.Y(scan_clk__L10_N1),
	.A(scan_clk__L9_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L10_I0 (
	.Y(scan_clk__L10_N0),
	.A(scan_clk__L9_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L9_I1 (
	.Y(scan_clk__L9_N1),
	.A(scan_clk__L8_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L9_I0 (
	.Y(scan_clk__L9_N0),
	.A(scan_clk__L8_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L8_I1 (
	.Y(scan_clk__L8_N1),
	.A(scan_clk__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L8_I0 (
	.Y(scan_clk__L8_N0),
	.A(scan_clk__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L7_I1 (
	.Y(scan_clk__L7_N1),
	.A(scan_clk__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L7_I0 (
	.Y(scan_clk__L7_N0),
	.A(scan_clk__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L6_I1 (
	.Y(scan_clk__L6_N1),
	.A(scan_clk__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk__L6_I0 (
	.Y(scan_clk__L6_N0),
	.A(scan_clk__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L5_I1 (
	.Y(scan_clk__L5_N1),
	.A(scan_clk__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX32M scan_clk__L5_I0 (
	.Y(scan_clk__L5_N0),
	.A(scan_clk__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M scan_clk__L4_I1 (
	.Y(scan_clk__L4_N1),
	.A(scan_clk__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L4_I0 (
	.Y(scan_clk__L4_N0),
	.A(scan_clk__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L3_I0 (
	.Y(scan_clk__L3_N0),
	.A(scan_clk__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk__L2_I0 (
	.Y(scan_clk__L2_N0),
	.A(scan_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L1_I0 (
	.Y(scan_clk__L1_N0),
	.A(scan_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I7 (
	.Y(O_CLK1__L5_N7),
	.A(O_CLK1__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I6 (
	.Y(O_CLK1__L5_N6),
	.A(O_CLK1__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I5 (
	.Y(O_CLK1__L5_N5),
	.A(O_CLK1__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I4 (
	.Y(O_CLK1__L5_N4),
	.A(O_CLK1__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I3 (
	.Y(O_CLK1__L5_N3),
	.A(O_CLK1__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I2 (
	.Y(O_CLK1__L5_N2),
	.A(O_CLK1__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I1 (
	.Y(O_CLK1__L5_N1),
	.A(O_CLK1__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L5_I0 (
	.Y(O_CLK1__L5_N0),
	.A(O_CLK1__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L4_I3 (
	.Y(O_CLK1__L4_N3),
	.A(O_CLK1__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L4_I2 (
	.Y(O_CLK1__L4_N2),
	.A(O_CLK1__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L4_I1 (
	.Y(O_CLK1__L4_N1),
	.A(O_CLK1__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L4_I0 (
	.Y(O_CLK1__L4_N0),
	.A(O_CLK1__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L3_I1 (
	.Y(O_CLK1__L3_N1),
	.A(O_CLK1__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L3_I0 (
	.Y(O_CLK1__L3_N0),
	.A(O_CLK1__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK1__L2_I0 (
	.Y(O_CLK1__L2_N0),
	.A(O_CLK1__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX14M O_CLK1__L1_I0 (
	.Y(O_CLK1__L1_N0),
	.A(O_CLK1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M ALU_CLK__L3_I0 (
	.Y(ALU_CLK__L3_N0),
	.A(ALU_CLK__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX14M ALU_CLK__L2_I0 (
	.Y(ALU_CLK__L2_N0),
	.A(ALU_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M ALU_CLK__L1_I0 (
	.Y(ALU_CLK__L1_N0),
	.A(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M O_CLK2__L13_I0 (
	.Y(O_CLK2__L13_N0),
	.A(O_CLK2__L12_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK2__L12_I0 (
	.Y(O_CLK2__L12_N0),
	.A(O_CLK2__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M O_CLK2__L11_I0 (
	.Y(O_CLK2__L11_N0),
	.A(O_CLK2__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M O_CLK2__L10_I0 (
	.Y(O_CLK2__L10_N0),
	.A(O_CLK2__L9_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L9_I0 (
	.Y(O_CLK2__L9_N0),
	.A(O_CLK2__L8_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L8_I0 (
	.Y(O_CLK2__L8_N0),
	.A(O_CLK2__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L7_I1 (
	.Y(O_CLK2__L7_N1),
	.A(O_CLK2__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M O_CLK2__L7_I0 (
	.Y(O_CLK2__L7_N0),
	.A(O_CLK2__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L6_I1 (
	.Y(O_CLK2__L6_N1),
	.A(O_CLK2__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK2__L6_I0 (
	.Y(O_CLK2__L6_N0),
	.A(O_CLK2__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M O_CLK2__L5_I0 (
	.Y(O_CLK2__L5_N0),
	.A(O_CLK2__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L4_I0 (
	.Y(O_CLK2__L4_N0),
	.A(O_CLK2__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L3_I0 (
	.Y(O_CLK2__L3_N0),
	.A(O_CLK2__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M O_CLK2__L2_I0 (
	.Y(O_CLK2__L2_N0),
	.A(O_CLK2__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX32M O_CLK2__L1_I0 (
	.Y(O_CLK2__L1_N0),
	.A(O_CLK2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M O_CLK3__L3_I3 (
	.Y(O_CLK3__L3_N3),
	.A(O_CLK3__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M O_CLK3__L3_I2 (
	.Y(O_CLK3__L3_N2),
	.A(O_CLK3__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M O_CLK3__L3_I1 (
	.Y(O_CLK3__L3_N1),
	.A(O_CLK3__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M O_CLK3__L3_I0 (
	.Y(O_CLK3__L3_N0),
	.A(O_CLK3__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK3__L2_I0 (
	.Y(O_CLK3__L2_N0),
	.A(O_CLK3__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX16M O_CLK3__L1_I0 (
	.Y(O_CLK3__L1_N0),
	.A(O_CLK3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M O_CLK4__L3_I1 (
	.Y(O_CLK4__L3_N1),
	.A(O_CLK4__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M O_CLK4__L3_I0 (
	.Y(O_CLK4__L3_N0),
	.A(O_CLK4__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M O_CLK4__L2_I0 (
	.Y(O_CLK4__L2_N0),
	.A(O_CLK4__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX20M O_CLK4__L1_I0 (
	.Y(O_CLK4__L1_N0),
	.A(O_CLK4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M FE_OFC3_O_RST2 (
	.Y(FE_OFN3_O_RST2),
	.A(FE_OFN0_O_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX6M FE_OFC2_O_RST2 (
	.Y(FE_OFN2_O_RST2),
	.A(FE_OFN0_O_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M FE_OFC0_O_RST2 (
	.Y(FE_OFN0_O_RST2),
	.A(O_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U5 (
	.Y(n4),
	.A(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U6 (
	.Y(n5),
	.A(Address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U7 (
	.Y(_1_net_),
	.B(n2),
	.A(GATE_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n1),
	.A(F_EMPTY), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U10 (
	.Y(n2),
	.A(test_mode), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U14 (
	.Y(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U15 (
	.Y(n26),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U16 (
	.Y(n27),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U17 (
	.Y(n50),
	.A(SE), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U18 (
	.Y(n28),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U19 (
	.Y(n29),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U20 (
	.Y(n30),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U21 (
	.Y(n31),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U22 (
	.Y(n32),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U23 (
	.Y(n33),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U24 (
	.Y(n34),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U25 (
	.Y(n35),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U26 (
	.Y(n36),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U27 (
	.Y(n37),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U28 (
	.Y(n38),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U29 (
	.Y(n39),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U30 (
	.Y(n40),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U31 (
	.Y(n41),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U32 (
	.Y(n42),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U33 (
	.Y(n43),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U34 (
	.Y(n44),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U35 (
	.Y(n45),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U36 (
	.Y(n46),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U37 (
	.Y(n47),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U38 (
	.Y(n48),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U39 (
	.Y(n49),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M U40 (
	.Y(n51),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U41 (
	.Y(n52),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U42 (
	.Y(n53),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U43 (
	.Y(n54),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U44 (
	.Y(n55),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_1 REF_CLK_MUX (
	.IN_0(REF_CLK__L2_N0),
	.IN_1(scan_clk__L12_N0),
	.SEL(n2),
	.OUT(O_CLK1), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_4 UART_CLK_MUX (
	.IN_0(UART_CLK__L2_N0),
	.IN_1(scan_clk__L2_N0),
	.SEL(n2),
	.OUT(O_CLK2), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_3 DIV_TX_MUX (
	.IN_0(TX_CLK),
	.IN_1(scan_clk__L14_N0),
	.SEL(n2),
	.OUT(O_CLK3), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_2 DIV_RX_MUX (
	.IN_0(RX_CLK),
	.IN_1(scan_clk__L14_N0),
	.SEL(n2),
	.OUT(O_CLK4), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_0 RST_MUX (
	.IN_0(RST_N),
	.IN_1(scan_rst),
	.SEL(n2),
	.OUT(O_RST1), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_6 GEN_RST1_MUX (
	.IN_0(SYNC_RST1),
	.IN_1(scan_rst),
	.SEL(n2),
	.OUT(O_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_5 GEN_RST2_MUX (
	.IN_0(SYNC_RST2),
	.IN_1(scan_rst),
	.SEL(n2),
	.OUT(O_RST3), 
	.VDD(VDD), 
	.VSS(VSS));
   RST_SYNC_test_1 U0_RST_SYNC1 (
	.RST(O_RST1),
	.CLK(O_CLK1__L5_N4),
	.SYNC_RST(SYNC_RST1),
	.test_si(SI[3]),
	.test_se(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   RST_SYNC_test_0 U1_RST_SYNC2 (
	.RST(O_RST1),
	.CLK(O_CLK2__L13_N0),
	.SYNC_RST(SYNC_RST2),
	.test_si(SYNC_RST1),
	.test_se(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   DATA_SYNC_BUS_WIDTH8_test_1 U2_DATA_SYNC (
	.unsync_bus({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.bus_enable(RX_VLD),
	.D_CLK(O_CLK1__L5_N0),
	.RST(FE_OFN2_O_RST2),
	.sync_bus({ RX_OUT_SYNC[7],
		RX_OUT_SYNC[6],
		RX_OUT_SYNC[5],
		RX_OUT_SYNC[4],
		RX_OUT_SYNC[3],
		RX_OUT_SYNC[2],
		RX_OUT_SYNC[1],
		RX_OUT_SYNC[0] }),
	.enable_pulse(RX_VLD_SYNC),
	.test_si(SYNC_RST2),
	.test_so(n23),
	.test_se(n26),
	.FE_OFN3_O_RST2(FE_OFN3_O_RST2),
	.O_CLK1__L5_N7(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   ASYNC_FIFO_DATA_WIDTH8_ADD_WIDTH4_test_1 U3_FIFO (
	.W_CLK(O_CLK1__L5_N4),
	.W_RST(O_RST2),
	.W_INC(WR_INC),
	.R_CLK(O_CLK3__L3_N0),
	.R_RST(O_RST3),
	.R_INC(RD_INC),
	.WR_DATA({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.FULL(FIFO_FULL),
	.RD_DATA({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.EMPTY(F_EMPTY),
	.test_si2(SI[2]),
	.test_si1(n23),
	.test_so2(n20),
	.test_so1(SO[3]),
	.test_se(n25),
	.FE_OFN2_O_RST2(FE_OFN2_O_RST2),
	.FE_OFN3_O_RST2(FE_OFN3_O_RST2),
	.O_CLK3__L3_N3(O_CLK3__L3_N3),
	.O_CLK1__L5_N5(O_CLK1__L5_N5),
	.O_CLK1__L5_N6(O_CLK1__L5_N6),
	.O_CLK1__L5_N7(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   PULSE_GEN_test_1 U4_PLSE_GEN1 (
	.CLK(O_CLK3__L3_N0),
	.RST(O_RST3),
	.LVL_SIG(BUSY),
	.PULSE_SIG(RD_INC),
	.test_si(n20),
	.test_so(n19),
	.test_se(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_width8_test_1 U6_CLK_DIV_TX (
	.i_ref_clk(O_CLK2),
	.i_rst_n(O_RST3),
	.i_clk_en(1'b1),
	.i_div_ratio({ div_ratio[7],
		div_ratio[6],
		div_ratio[5],
		div_ratio[4],
		div_ratio[3],
		div_ratio[2],
		div_ratio[1],
		div_ratio[0] }),
	.o_div_clk(TX_CLK),
	.test_si(n19),
	.test_so(n18),
	.test_se(n35),
	.O_CLK2__L13_N0(O_CLK2__L13_N0),
	.O_CLK2__L7_N0(O_CLK2__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   Pres_MUX_WIDTH4_PRE_WD6 U7_PRE_MUX (
	.Prescale({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2] }),
	.div_ratio({ Pre_div[3],
		Pre_div[2],
		Pre_div[1],
		Pre_div[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_width4_test_1 U8_CLK_DIV_RX (
	.i_ref_clk(O_CLK2),
	.i_rst_n(O_RST3),
	.i_clk_en(1'b1),
	.i_div_ratio({ Pre_div[3],
		Pre_div[2],
		Pre_div[1],
		Pre_div[0] }),
	.o_div_clk(RX_CLK),
	.test_si(n18),
	.test_so(n17),
	.test_se(n43),
	.O_CLK2__L13_N0(O_CLK2__L13_N0),
	.O_CLK2__L7_N0(O_CLK2__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_DATA_WIDTH8_test_1 U9_UART_TOP (
	.RST(O_RST3),
	.TX_CLK(O_CLK3__L3_N1),
	.RX_CLK(O_CLK4__L3_N0),
	.RX_IN_S(UART_RX_IN),
	.RX_OUT_P({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.RX_OUT_V(RX_VLD),
	.TX_IN_P({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.TX_IN_V(n1),
	.TX_OUT_S(UART_TX_O),
	.TX_OUT_V(BUSY),
	.Prescale({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2] }),
	.parity_enable(UART_CONFIG[0]),
	.parity_type(UART_CONFIG[1]),
	.parity_error(parity_error),
	.framing_error(framing_error),
	.test_si2(SI[1]),
	.test_si1(n17),
	.test_so2(n14),
	.test_so1(SO[2]),
	.test_se(n26),
	.O_CLK4__L3_N1(O_CLK4__L3_N1),
	.O_CLK3__L3_N2(O_CLK3__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SYSTEM_CTRL_BYTE8_test_1 U10_SYS_CTRL (
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }),
	.ALU_OUT_VLD(ALU_OUT_VLD),
	.RX_P_DATA({ RX_OUT_SYNC[7],
		RX_OUT_SYNC[6],
		RX_OUT_SYNC[5],
		RX_OUT_SYNC[4],
		RX_OUT_SYNC[3],
		RX_OUT_SYNC[2],
		RX_OUT_SYNC[1],
		RX_OUT_SYNC[0] }),
	.RX_D_VLD(RX_VLD_SYNC),
	.FIFO_FULL(FIFO_FULL),
	.RdData({ Rd_D[7],
		Rd_D[6],
		Rd_D[5],
		Rd_D[4],
		Rd_D[3],
		Rd_D[2],
		Rd_D[1],
		Rd_D[0] }),
	.RdData_Valid(RD_D_VLD),
	.CLK(O_CLK1__L5_N0),
	.RST(FE_OFN2_O_RST2),
	.ALU_EN(ALU_EN),
	.ALU_FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }),
	.CLK_EN(GATE_EN),
	.Address({ Address[3],
		Address[2],
		Address[1],
		Address[0] }),
	.WrEn(WrEn),
	.RdEn(RdEn),
	.WrData({ Wr_D[7],
		Wr_D[6],
		Wr_D[5],
		Wr_D[4],
		Wr_D[3],
		Wr_D[2],
		Wr_D[1],
		Wr_D[0] }),
	.TX_P_Data({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.TX_D_VLD(WR_INC),
	.test_si(n14),
	.test_so(n13),
	.test_se(n44),
	.FE_OFN3_O_RST2(FE_OFN3_O_RST2),
	.O_CLK1__L5_N7(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   Reg_File_ADD_WIDTH4_RdWr_WIDTH8_RegF_DEPTH16_test_1 U11_REG_FILE (
	.RdEn(RdEn),
	.WrEn(WrEn),
	.CLK(O_CLK1__L5_N0),
	.RST(O_RST2),
	.ADDRESS({ Address[3],
		Address[2],
		n5,
		n4 }),
	.Wr_DATA({ Wr_D[7],
		Wr_D[6],
		Wr_D[5],
		Wr_D[4],
		Wr_D[3],
		Wr_D[2],
		Wr_D[1],
		Wr_D[0] }),
	.Rd_DATA({ Rd_D[7],
		Rd_D[6],
		Rd_D[5],
		Rd_D[4],
		Rd_D[3],
		Rd_D[2],
		Rd_D[1],
		Rd_D[0] }),
	.Rd_DATA_VLD(RD_D_VLD),
	.REG0({ Op_A[7],
		Op_A[6],
		Op_A[5],
		Op_A[4],
		Op_A[3],
		Op_A[2],
		Op_A[1],
		Op_A[0] }),
	.REG1({ Op_B[7],
		Op_B[6],
		Op_B[5],
		Op_B[4],
		Op_B[3],
		Op_B[2],
		Op_B[1],
		Op_B[0] }),
	.REG2({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2],
		UART_CONFIG[1],
		UART_CONFIG[0] }),
	.REG3({ div_ratio[7],
		div_ratio[6],
		div_ratio[5],
		div_ratio[4],
		div_ratio[3],
		div_ratio[2],
		div_ratio[1],
		div_ratio[0] }),
	.test_si2(SI[0]),
	.test_si1(n13),
	.test_so1(SO[1]),
	.test_se(SE),
	.FE_OFN0_O_RST2(FE_OFN0_O_RST2),
	.FE_OFN2_O_RST2(FE_OFN2_O_RST2),
	.FE_OFN3_O_RST2(FE_OFN3_O_RST2),
	.O_CLK1__L5_N1(O_CLK1__L5_N1),
	.O_CLK1__L5_N2(O_CLK1__L5_N2),
	.O_CLK1__L5_N3(O_CLK1__L5_N3),
	.O_CLK1__L5_N4(O_CLK1__L5_N4),
	.O_CLK1__L5_N5(O_CLK1__L5_N5),
	.O_CLK1__L5_N7(O_CLK1__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OUT_WD16_DATA_WD8_FUN_WD4_test_1 U12_ALU (
	.A({ Op_A[7],
		Op_A[6],
		Op_A[5],
		Op_A[4],
		Op_A[3],
		Op_A[2],
		Op_A[1],
		Op_A[0] }),
	.B({ Op_B[7],
		Op_B[6],
		Op_B[5],
		Op_B[4],
		Op_B[3],
		Op_B[2],
		Op_B[1],
		Op_B[0] }),
	.ALU_FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }),
	.CLK(ALU_CLK__L3_N0),
	.RST(FE_OFN2_O_RST2),
	.ENABLE(ALU_EN),
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }),
	.OUT_VALID(ALU_OUT_VLD),
	.test_si(Rd_D[7]),
	.test_se(n46),
	.FE_OFN3_O_RST2(FE_OFN3_O_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_GATE U13_CLK_GATE (
	.CLK_EN(_1_net_),
	.CLK(O_CLK1),
	.GATED_CLK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

